PK   ��X��OZ%  j    cirkitFile.json�]�o�8��W�=��/�̷y��w�Ә9�~�n�DM|붳�ҏm��~���-�v�������*���UŢ�e�0�l\�v��.���lpK�ppg�G��i:�Of�z>�}a���_��I���&����|fg�8e"eF�Dڂ%<�l��R$E*������q:�}�nx���:Ž�p�s�z��9U�4�L�66�°$�2KT�2[��R����6��҈2+�BH�pcub)��k.󴬬��]��#5����Z�UElN�Tg2�UI�g,�e�x������
ѲĴ�1-+�4rza�'r~�J�a����9r����~p�@��D�|!�	C����!�����jy�m��Q3��aP�(�N��)�m�j��:#�i["�\4�i�,aH���˱&� ��KS��V��D&��V	fJc��Y?0!��ZF���,�곶���,��P�Ėi�#I�O�B�Z���6�0-�\|Pˡ��(s���VZzU�J���v�����d4�p}-����a&he4�o��s��,�׉��2�;���
- ���rh� N*Dˡ�hH-����a�z�A�M�	��x�Q�A
��{�iehhŇ�x��C"��ô�Z�Hh�C��@۰������OD�$h�a�!f�5�i��R!��`�L�(�2�����OoX�rМ�rb����L ����i:���N�^g�@��]-P(B9�#�l`���!}�'ؤ "js���vW��O����Oi���A7�"p�Q��(\��RU)�%���\2�J�#�dQz$W\dVU.*�,:�"�7zI_�\�L1l��L�0lx�N�8l�@�46RH�b�$�i��J�c�6�UU�t�]"o?3�	�M�b���-�M�b^�ܠƦA��i�P��8
oP��Π�ŕU8ܰ8(fGm1t��)*�r0�Э��d2P�ܖ8,t�!�,t��G��?�#h*��?M�G�,����kh�;��k8��ѵ	��>�6�ԇ�&p����N^����k4�{8�&f�i���	�.=�JB3���4�y�� 3�Gt�.M�����
4�w8r����*`/���4�w�4��f@��9�:@sn�{͟m{��[֦��\��>�3E���\h.,
����%��EFᢢp�qP	�q�K�����/�`�$�I�8 &qPL㠘F��qPL㠘�A1��b�4�i�8(fqP̎���s9*8��G�����s9:���0<����s9:�������8�=�a�sa���q�;���s9�nh.�娲��0<���ͅ�đ帎��0<�����s9>����\��0<��x���\ve�:t�~�WUa�I�ipK�p�q�������Of�������D1r��u2�ޡ�Fm�r\���/�)�Y��HM!e��*u��"Q��$e�n c�,�����q��PȠ�
��.�j�c��3(dPYLۡ��IN�)�c�i9��>��9u���Z�-�d�i\q0�eLA\xZ�<TT.�4ƈb�g��vVNN�a61-c@��ZF����	��0�_L��__p��qe��><Q��Em�WTa����it(�����~~�-�l	0\�l�=;��G�1f������!�K��ۊAP�ː�"�{��c(� �?}R��bR��D���?`�
Z��ٌ}~M?}��|���K���&�C2藳?�Ѿ^�����g>����[v�e#��K4��5.3R��g���$����;)���C�۵�ȇ�۔A-���[�ͬ�+�z�t�Q����e�;�D�ndF��S �]�ƫ!C���42�G��/z��E@O;��iw�
_��0��"�"`k#�����E@V&F�^ �^ �>�a.Q��� ��@���`�9x	�i��99��Y|�_"�(>
� / ��� �(�ţ Y�4I��=j�.Q�W�H��T��*�D�0^����a ��?l	/QA�� �8S6�1�7�򴧱`;cb,���C~����h)�=��ۀ#H�ٺ�Fl�@�1�	d	��!��,��K�,�z:��Z�'v���4^�E��J�8�tl."Cp0�X.�Ţ��i��s ��6��G �3w�d�T ۙ;_�X�1�6�vN/�%���,@xu\}{�����O�}�#� F��cO�^��,N�����ΎV�|#ug�ç/EG��$�Pl�
�|�B�(c����,V��e��a,|���H�ӫ��g;��Y�W�(`ex#�2���4��c����vj�]�����\�����h1���B��O�B<�A>���I���U�b�������~���p�/��K�/~7�E�0�mo���=��{�ä�^�=�xr��)�}�|��ڕ�������K�:�B��wi:�09n�{���X�6WB��9������PsI$��� �2肖
�a���%X�R,l���[�u@���3Ĵ��4P��Q�@ ci��Fm=w�4nYb�:��@}�N1
e��n��-��}�U�-v�s=҅"���-v���;�9�c�)H�ڊ����;�f{�P�z�w`�/�Ƽ`)�_��b _
�w|����O�/�n���ݚʨJj�R���/d���؅��f�;���?�\�]���B�6����0�=3��,�>�;\�4�0�b�RЫ�CVz�8��1�b����+�[�X��w����Y�K�[��|�x��_��G6��'���B��훁����U?��t��q�����f���,
�%ofi3��1o�E�ƒ6���Z���� 6�oP�Fs��7������\l�5f�K��Q|�d]��_�&��w���X�������9F����2�;/8D>��8�����=tl:н��w��qӲ_���Ř�nGh�#���d�s���.J�0�ƭ�!F{�Y7�E�����#��ޅ� 1 F_�֍?1�oL놯qЗ�u�_�8�{պ�3F�Uk��#���n��Xpq�&�0�ӑвr����0!�y�©�4!�y�"��4!�y�j��4A�y��`��%�4�
��x�������vڄ��#�S��Mc����Y�}D׏h��p�>��G������=f�GY��\?��Gj�Hu��#�yD6�A��A�}�v�l��tǊlzM��&��"��"�~�n�ɦ��s��9�v�l�N�}����_��t:޹�d2����dY{���4a阎�g�`Ǌ����,?�7�y�vR3�M�-_��^/��vQOl��y?�����_֋��w׳�y���O��f����\y�<�&����my7�����tp[��Һ�K��m���S��la��0Y�rp[�޸�yof�)ꇅ�{)��.٣�e?/kױ�8Y���I=��Qx�PNGLũX�T!Fԅd4]���zy_9[�*/J��\V	͘2�}J����H���b�����bٴE���lY�Y�bʋ���q1+y ��dQL�Z�oIGbH�w���	az$����k��K��Կ��d��i@Fl�t_pr"NR�G�gJ��G4{���ap��G���8QR�5O٬���w.�X<L�W�����:2��̈́��
����b�|�=��%�ie�D�z�'�sI�B[�U���P&������f(i
SƭQ�T�jެH��'|��O�y��6J�����<��O ���ή��@k֌�q�	%6F}:���ɤL��l���y�U�SV2�l�A��i@�Ir��(����O�7E��4�K�]���#�hJ��6�CgVɈH�&��*KOH������ !I�9_�#)���R�P��G�3:�[�T� K}�Y{M���Rg�F�,��tٺ���)e��a[J�e~:2?���"�ξP�C��c���/��u�=��1ήٹyOe�	���A�0�l��A���ɽb��j�A�U��A7gk�M�כ���+��C�� ��/��R���4�d��l9��MY���&�v�]o�)�<X���9)g��f��	9�R��h{6=��דn/�O��ܸV"QL��h���f�!{��q]L~��,Ϥ�(�J���Ʈmgw/!�{�*DG��^:�fw�����k���L���6K��ȏz!�Ԓ�U"Jm� 2弫�L�*��nr��w�;L/L7�=�=��'nY�����o����E�Vt~E\t���~隱�qk>�jMOw?r��]���9���q��n!##�������>)+s�S�H��D�HLJ�D�����s
�'�����B[��lB
|��o��[rߙd<@���O�Z�)�	j��r;t<Ћf����f5�t֭� v�.C�P���s ��ڎ�d@B�HS�$�z�~ƀ�P�$c-U�ڟ�!:��� !�mL��fP�]�; �k#X�a�}�MF��&]:����.�_�6������`�O[wo÷�I�|R��W��P��	�$K��lRT��.l�6����t�֍���O_���,�v��,T©uFۤ*�y��<��e�o罂9��f	�έs�]%y�ܒ��L��V��{�f����R�db	!�	,2�rY:�q�x��lѪ��W�_�g����%�'?�M��g��d�҉"�N�s���,)3�KK����P�`�y���p�rQ��lɨ�����HT:%�ȕ�=\~�ΗvWᚤ��Ie��K&�$��P"���G^���ͬ��=�
�����{.�W>k8�?�5��y��.��7(�}�z���+˅].�ϾɐS>�&S���d�z0�:��L���fn<ቭ$�q}*0����Ĺ.�2q�uaVJ�*���} ˋ�Ry�9j̔��,7$���2'T�����aN�r�F��/������>B��a��?�>�'��������/o��nn��������b���S��م������f�<�[G������a4�����7�Y���������.���ک-�-d���`e<���/�n;q;�̛��|*v�[����Y�x���9�����hj����}�	)����>N���I�QJW^��m�	�7MՈ�T��O�W?���Eস���۝��[ן�؏�p����x~�slT��Uo��r>�~=��rv�
�� +XYl�ja>�S4��񤻟Of�kS�5�j������k���&4Y�Oo���ﻮcBw#gO0��T�U�j�R=Ż���98!��T�
2N��H�b�1�)@�0*�ΝG��꜀t�؏�s��	��t������2�*��eU�0a���tI�<A�X�$g�ro#�o�����BB:�!i='�jv�"��>A�'��j����=�qk��Q�����������_�:�rMc*f�a�_"+l�O��d��mQP|�.�uߡ��x��x��NP<\�X���Q|�7?>�;d{�[�m�	�Ű�cX�."k=�tgi}[eup�wȶ�(�A�w�B1�̪*f�.�i�G��eT����t}0ZoQ�ޘl��	D�ڔ0:n�F4���ᢹ}g�}�H�?�z�!ӻPy����K�@�Sau�hTU�E�,H�p,x�|��C*<Zd4�50�?rU�YN�E�G�0eq�qV�o�8�پO�%�x�����J��F����N�q�����MF;���l[�+N�<7q}'D"�g�"��!ax�Ț��.٦���D����#��"9!=q�p��qV�b�"(��~�c��)��N#{)�eL� WзDD�|m�Kw�c
����~�s�x��:� }�Հ���h�#�J�cY���)V�<&2���X"#�o��;
�kS��G�� N����)cUL``$�n��� �@.މ��/�A�M�}���S���PU%��d�o&���9O���;)�j����F�g�N��B���7Q#X�T}kTlh�wU�❺����W�����p<��mTV��\���=y����E�0��6Y���?�zyYDޑ�*<�'�UTx�WA-a�Y`Ӥ囀��� &����O�����.�1��ɿm���=������j��6y�Σ�~1�_[�?�e��ܯOm�_�PK   ��X�<1	}�  � /   images/02d8db12-ba28-4e49-8e56-db179b980a39.pngԼ�WSY�>�Agl�b�HDz� �H�)�AJBI(c���@��H��B��!TC'�J(��N|�x���keapg�{�庮{�s��=��t^]M�!t�
���)�/�]�ׯ��~~P�Y� ��f�q~��N|�7��x�S屧��SO�'�6 ///a{G�'�l�]�m߭�_���+�5�N^��IN�IY��t�MQ�&���w߻h����wU��p��]���x
o�qOֳUm��C����Iw�M�����_�Fkp�7JQ�:o�V��o�o`��Z��dW#8�Pv�F���*#蟟4��G�cB��ܯ�������?�}���~����;ƺ�N�M�!Pu���%��cS	�=�zl�8�co۟?�;�����\�$�����;|gGo�m�'�ODۏr젩!!�e��H�P3����w�f]����E�k�p{�� �����-7�������� R~	<�����0��,T_�ӑc �r[�k=�[W��uEO�_�]+	}:�պ:zE}=Uo�[�b�5K<�Z�����V�UU�o�zE�<�]f�oQ�.Q�}
�����;�Ue->�\����D]����-��.��I�յ~b�2+��)2�32+wV'�B�kY�@ A��+��⡃A�z�66�L�������;m��ѣ�7�$��]��R�^Q�=�svgn~U�b[��oI�ԉ���x�O��Mr��T߀rR��P�����o񯣼��NbLMYߍ����+�u��G��5�I,�;՚I[�]˯��zXӋ�M*}z���������C��H*s��J�ҳ�k9{%(+��c���_�xu�K�@>iY�����وG��AF���L�Oo�f�q+�T�y<7iX��֣	�6\���o�`Q�F
̆��p�a(c|+|�{َVG�����2����a'�g	p�-��+��=�D��V��(AGN��d<N�#1�v���s-��u)_���	���`"�
��qj7�'4��m[a�,ӰQ�n�<G�ؕ�_�nLI�
��LB��fM��0�W�]ܺ2�H�i[�cSg_p�k8������^���^ٝ�V��L0#H��^>V�GQB����s:�ɺ"=��PV�Nv7q�\�pEE���
%)��f���}�_��~����	K�s;xz]�V�3R��E�`I�@▝ܬ�P����4��uXKV��.�>��4}��S���;�z@�ަ6���ҕIUH,�	����	 ���
�C�%�k�9�Q5�w�.�����V�s��3ݑY�*-ߊ�'Aaw  H�e��	:�Џ֋*Su����L��_R�S!��0�_��z!z�Ŗn��DfŊ�㹵C����	�0���]�Թ�.�r��Κ��!��������[�6���s�KvQI6����z�O��n�i(��$��(����z(�jC�5�_�;R�b�y������Z���{����՗
e�Sw�ν�2�����UZ����_�2?ɤ�/��럺�S�}�/�3���[GL�|��7����֕�TDrX\�J��Ҁ����]����Y�@~�GzGD� ]�G��*u��E7aa�2\g�����V�H$
�/�<���B���`�?Fo
���Dxi��)c��4K�=9d~f�%ں� �;v���9	�<����Uj�(���y@�N����ގ��	
TJ?Z��/�H�so��@ܸc�Բ���	M�!��eW��E��h,$������nz�n�9r�:;���T��EOP,N6IGZ�+����;��c��Q�h`ߞ��Xݙ��rQ`i��*I��r�b��[7�7�G4t�7ǢR:hrͨ�����c�jd�Wa�3�vo���Ɲ��K�&~�$�'̩aBmN�(�<�2��l�����]�#�|7Q�{%`g0��C`1&�eT�i*&b©����Ӡ���:`7=iN��ۻ"=�_�`�U�3&����O�����95u���8�NY��%�kq�����+>3P.L���E���1{~�u���&�*�4K���D�ku1f��k=���
�y�XvD��
c��:���!��" g-ѡ�J��~̜�3���f�����A��z��w�#���L��,���:'I���xn�,���Bj����U
����Ӊ��T��2�L�۱���T�ʾ>���˱��4�vnw'���UK����}��wc�i�:��u\��-�3(�`'�us��>���t,�H1-�W��u�TF{oB���l�P��Α���6l+����^�.��vZB�IO|�((MG���BB�	�iȃ�\���ݏAPװ]�U-�S��#�tg����.�����i�O�!�[�>H������k�&6_�ᓀpf�.dP�aQ���}ڿ���9����kO@'�s�|�����-=�
�q���qt/'�"W����ǫUk�m�?&��z"P����N�����Y�~ϫ��������I�o��\���/��:�և��DOqyӟ�9�M�o����?������z>�Z9�?��}%RW�;&<`z�L�Ag��"V���O�,9	'h�3�� Y��s�F�e��><v�W5�z�} ��/����~��O�nI��Du+T���Y'��D�����%��9��T�OM�c��K�랦O���@Q�Ձsk��2�i׺}K��^������OW�� �ZG}qy_��_�eL�\��Mm �q��%��<j�3�'h	=P:����Cos,D9j嚶Ю0�r�6���dz�ŝ?6��T���#0�����O":�?��NS. 7/�r�Xx�'� �I��cT�VFH�HD�[��Y�� �`6�$�a�1G�+�����Ma%�
 ����i~�x��z�q�~t/���Dvѧ"މ_WE_f�EG\�VU�oeu��Q'����P4��:�^캵:R�h�2^q����n�)dԜU��M������7��\�7C &�EՉ��)yJ��{�૜��Pn��$Z��K齷V�_������zC.����Ma���mb=�}��������+��2���zr�sC��0�]��xq�h�:RSY�v�u�u3�]7�4$1��M-1}�:����s!3:2�Y)n�%o:88j����W%m4�d�6���INM��d�?!�{7�߲�Ȝw���E*�0XK��GmeZ������f,�}��S����D�G��]��K���C�3O�*�(C䮇ϲ�<�A�h���.����]���R�XB�e��g�^f/j�/��ㆄ��odޚ�������H���0�_���� i�3�/��e��sTDK��;V��D­�o�����Ab��U�����Fy�ԋ�i�&#�����m������%,��{�4/\8���7��"ʀ��Dh�	g�0t��}P(rJ�`,�+6��e���U�:��@ϡ�r7p�k�1o�n����� 	������n.��]E��Y�dT��D��±�vH��٣JҘ����j�@Y�|� 1ޜ�H�z�b�$�J�$�� =J���N�"K,ZQ�$0q�s��{�E���YH)���i�VI����o.�_26���B_�m[���jy�{fJD��&_�(L��4���\=�e�-����q�`9�F���HsT%I�//�G� �����ط�)B6Ϯ�}�񵄭�/\��+�����V��U�5�gd*������k%�>�����3_�r/u�(�HA�'R��-8��=��z+��Ο�B�;~{��Q<Q3Odl`��徃
}���g��l8�Aܬ�N��Կ[�`��!L�-�kv���v�1�|����\���c�������
h���=M ����� �ӯ� ���M`-B�^]�ˈT���J[�����3����d�nJ"��&�7��8����hvu�%c+E��+�~=ېŝ���I��
�|r[���Tw��$?���e�1�e��U�q7{蒄�vD���6;���rī�' ��W=*ζ�1�X!�Tw���e�YB}eg�|���2�j��d�%��S5�C?�P�gK�K6�7�x��|�>?<�S]��ƕ#�_0ђd��٪�!�_>ǎ��\?'W9~���c����;��ذ�ig��@Ná�Аr��/i�ZLl(����S���=�uȿ��1(F��i��UQ�]��H�7�b�qzt�4ݗ�^f���%'|@  ׏��y��l䷬��.��X���s�e~���]sښS (󺹪^X�#�� Ҍ����c�f���\ȯ�z����QQ�n����$G���Dz�59��>9s�]s��kv�L,��+̙FК�O���_�-� 
L[��]����9P��S*u�;,�D���g�3���v;�ɂ��D�������`�H}��B�Il�+�����7�j*����+��4�Yř��4�o~4`r>`���V �~���F��52�K���#>�sWUb��"����lٴ�|!�sF�.���[JB�'�u���nd�E'Q �\���J`x=���;ueܠ;mG��-�ry� *�I���v��<;��B�H�0;�!^)�2Fn���#/Fb�kfj��`��MطT'%`4 �%�kJ��ӝqZo��Z��0��rJ7�|SC�}!1��L?n���j����0g�N�z����  m�@Oh�	��q���HEw�����)����Ήa�ȓB��U�Q��Q��@���_i��)"�*�v�o[�M>.�׹aV+���!���W&Gb��Q7�	�Q֢����<�v��{m:�����ݕ���T��� ����78����b�;��-����a�X��74�>0����@c&Dh�6�9[�ʥH�D~�#1�G��E$��uӌ�ë�Eb��r�P�܂���Y簤�9�L��a����5�[7r��e+ٝt�	�&�͖I�_G'�J �q�!�u�D!]�%H���� ^n?ʟ�埨�D�#ߟt8�Գ�}0���T�inA�V���L��@GhFA�G;�b��d9~^\�]��KY�n�����jR�! 3Lr
ө��CXLX�$bb%}e�	Xuko|��]7�[�;Z�@J�)0�@�B#X
"B�\�!>��wv��,�+�
 +��{���[��>6�I"S8�D
C ;m�K�+u�J��נO��d����͢�I��.��P��^��?*뽞>`85#!��
�}��lEB##D_,�����|(�p��wQީd^g3Z�}�՗6f5=�پeq=�с�ST#$�~9%SF�e�j��6�V��I����hNQM��<���g��j�m�W� "fWi���M7�@/���F}����'�'�5��y���z���6'yl�#_֑h�1��Q�[ݫ��kp�a��K��4ٷ䰋u�
5k%�!"b�~n���)����`bb��P��������^j<�{^:c��*�V�B��A�p�����r�YZRؓ;pɃ��"6���G2 �W���2^�����zڊQ���l��<��X�d%h���H/�h�gUH��Y��>\� ��mCֽ� ��ҭ�-���p�W��d��p���O��N?��c���%~F# `b3Qg�����g�ʺ�<#�_��Xb�:�9��'�W�~�j�Q٨iJ��>̻)�Q₧kh1�: CXm��!�K��25�n��(+m���eGE��Llb���؅�ͱ/�nl�нx�6������I4��\	9������J^j9B ҙ���ތS��/�L�I,Ln�O��Nٻ}�JQ�I����7�H-��R����籓���Z�B�U�\�y^�z�t�������ˀ��!�M7��H���S$	��a��@G"d��=X'�+�]/(��\O���r�u�_N��c>�����΀��(l��9����4z>����xZ;����d]�fv$䢔��BQ��K�W	��`��g^r]Xz���PXN{]"���T��!2Z/��AJ���C8F�Vrn�KH�����ٖ��,Ռu��ŏ���M�Tf=�ԟ`jN��Bm���t����|����p�R=¶ni,*��Z��@#']��0���:O�Ά��Y5l�m��i3��Y	U^qp	����h�/��6�,Z����:CW~��BF��]0�.�?)�2���r�[��9�ԡH҈nLy�����V�d����ӌh+mE�JBY�2b8�^]����/w:��U��4v=�f.��Ѵ��	���k�lV�(��[�)�8��	���ڏ�<׽sX��-�2�C$�U�'VN#��s�o��<���*�����㏧��nݮ���޸|Fl����ܽ�wz�+ݞ.4���cv�z��^G/IGم�Z]ь�YPe���v�[��r?y����*�a21�����	��}�u�uQͻ�А?�+_Xs�ͯM�#/깩Y9W	t�n��/�;�XԊ�ZԖ�Р��Be�HBnv�=,e�
t����M�~v:�����`V�H��
�I�2��v?%dmu�D���O[��ɐs�
�5�d]�U��;ŕ�9���^J!4�K�k�Z�ix�n��#ũ��|�^ڐ)R�Y���K���L��>6�L��� (t<���@(�r]wA�~�&OgWB�&�/��FAN���0���O�����b�tlNx�e@�h&^�����I4 s2Y��S�4�,�h�`�����m�yU>����F�
��	^������s�I����:a��~m=D�	Gn�R��e����Ӗ3��=S=v@��:�zm�Mї�v+�������>�-��h�TU����}q�C�2���c._f�ҏ8lT�C4��bT^���⿼gi}�E����܄��̴��:[�	�H��s��-m�Y����fJff��UvQ��\^86��-����l���V��`�F��0�����`���ª9���>�N�1B8�_?T<\�^�d�س��z�MS�J�lJ�C�{
��ukK�d^)�+{�FϹ���*[��ŝr6IS:[����,̪ �Vy3j�]:����a�,��pp=
�����L�ſ��ϣg���35} �z9%z�@GN�s�޵Վ}u�聄����|\	�����P���Lβ�(.S��=�L�yX��a��1z��6�>� ��>����S�Oت�\3F-}rR��V�Ji��xrB����y���n�Aq�j�l~��|��b@6pQ�fc���vJo��\Hs:D��zI�Bq�@������\=p�멃���L@i�oma3"����	�����>���PtxԞ��΃��h�ө�n}P�D�\�t,�i��w��]mA�D��7>���)G�N�~y�n0���K�"�V�p`�p���k/��~za#�ޅ�~SI(���+HY�s���\V̗}
� �8w���zs��g�`��Ԝ�v���.�⛫&UE�>��8!��}��m������¨B�imr��S�*1$d�{e�s�c���r*-V�$��Y�ܧ�8��򪬏���7�	�o��E�H{,H����zF)�c�r�{��*�R�<�^Z������/� P�>���Gmj��˦��Fքm���;�{a��
l���5�BY��I�h��4~xr��	��w�$C3 .�ອ�-L�ظ[.m��=80�"j@���[P�� �K�X�&m�v
��мV�<��M�����(�T��c`�l% n �_z%��G��������e'�I�V���qC��s��l`�df���7��n[����I��#���B>�s$�_�s��3�	�O��{2�(L�hgث7��$@JC��9~��QC�/gb��υb��:\��q���U��}GhQsW�B�sZLd�LhB% ��"~�7x[��Q�
*�\��Z��q���ؕ~Ӡ(�.~���ڮ�zC����1���t㨔�8_��r'��[1���{�c)�f?����g4�ۻp�n���-m׀��4��[�iCO�L�����a|��%��b��������On��;ӣ�7�p�Ϸ�c�D���
b{�	���2me+�@�ɒ�o�yG��}��j�b�4�vx���ƍ|��łi��%���N8E���]�ɭ��[:*VH��#��z�����=��lrIxٔ\��R���T|�ʲ��{��?Q0��D����3�g����!^:'�N��:����-O��� ���5ӱ�%nȧ���y�-+���+�"�qˎ%�o��ޏ9J��Ig��D���r�!�J6�p7�㺥����37��ĩ���������^.��,hC��Vy���pk6�D� �7V��N���U��`��3b�$�,�w]o���Ww8�v�\?�B!ٝ��<���r^֧�і�E�^^
ۂ�=�!�~���[΅1��G���Pw�p���Q�+;M�ML�"�:t#}��ـ��*��ǎÿE��89���'�L�ï�}�|7C������0QgT���)�ʪ���-�~�p�z�?��J����t.h߸��V��J�j�=���>�e��ב)�WZ[��ʼ1"g����y5������ZZ@aa��;zUo��/��S�3�0�������.��Rw��u�q���R�c@N��i�?��9!�)-�H�J�Wt(������gE��Q֣�+l\+��txP�i2��!���'���q��/g3�����T���zl����z�ab�f�����%���xT��|��6�;���JGs���$�#W��L��/R��/e��4���
�����?b����� P��Q#��Zc,DxQ������Yv���;�R�{�u�} ���՘ͻ�᪅��Ċ�}F�� U[O��*@D~+�П�����[�SQ��ʋCsE]�Q���@��Ǯ��/��x2���Y��e���X�L*n��}B@
�:����l8�m0���B�-F�:_�D�E�t<kBN���tRN���S
H��CBI�ľ�����v�����u=�l�3�iص
q+�1f���z�h�"�Ql�,���g���h�vh����_fqi� A���2'�t�w��
���I׷��܆��F�P��Qte5����;��nUT���cs���ڼg����t���T}o_rە�Do�&�'�r�������vK��d��FNDʕ��ˇ�%JJ����=�w.�;��X!�?1�9�v8S�b�57̐Y���/s��*�ސ�J �<�[���`Z������T�����+�3�[��֕�_�a�-��!��Z�;H��p�^��y�V�]N���w߭�}�ķ��]v1Y�M>�et���n��e�-⥿mG�y{�@	��拾'@*^�F������\۟�Y�|�G��{�C��BK��M��WM`~?w�ki3헙e�׷:W�z���B��sD��Z�!�	��mj���V�|�J�k�c*���
l8���B��9�cTV�öRt�����9G�����*�f��l�0⫁�e:�[<|QWG�6����@�)��jҵ�7�"Mp�Ut�n�e�+H�""җs>2���~����%2�_�=��tV�/@&u��9��ҹ�8����6�VX4�ڶ�&m"��P�����-�~����uB	�Zr�p��s	�%��_�#�?���|�8'��U���b����2��UF�7kk�/�D27_n������z�=̰H��������w[��B�������S����.J�M;�p<���rtj�v��2�I��I��+�;Ӷ�5�/ِ�Ľ�g�TF�����v$��>}n`rYv=�(�y���-[��u�w���i������NU��G�@�G��~��1�NyQ`}��dAu�,�D��d޷ E�J�*V�I���$�ń����hSmVT��N�Ƣ���M�U֨��������Y'�R���A�@��K���7� 	>f���B���69�(�aK����-�I����)ϫ����bX<���宥Z�����������E�^��K����Z�%�1�<h�ښ����42q5�B�i�D�ܤfm�sw �����oo���*�@��\�)� �/H�����pI���̇�6�(EHOW
�m�N�=4�ND،�fW� ��4�%�с��)�Q�Ý%�N�����*[��t��y�6?�/�!�r���tPX��*�*�S��ޕv��Xe���>�e����m�?[�\��s��8L�SZ��^��V��T��aJ!�C\���
lm�;��=Aa��W ~g�	�9B$���%6��!zغY�U�n c1Sȝ��̺��>���I�V�2�+�&�"��?����)3��)l}���Z��χ���͊X�D����I1Z*��;�5���\@�T��,X�e�UE
�izxȋ!x�0aLa��t/��>�Xz�e�)�-E�_tx�~���4�%Wc�]Rp@g� ���(�Eb�o��`��:?�[
 [	�e@oʺ�h��Dۿa�m�N`�������?�~qm�5��Y�D�_���E��;3�4���N�ڹ��x:�ʚ����|º� %����������7m�e� ���5"�n-_�(yK��W�W��9G�
U�R�|6����T�ls�����"�(3���-��h��vIN�d�XtX"�K
b
LDH���K5��pn{.����Ão%�OV��)�[w[���yAv&q3�'٬�w{t�̞5���� ���[����Ȫ>�y"�׻h��t�'��.0IW ���D1NE�,�(1ʼ�����-sF)����p����FzD]�LV���|>�4�jI�f�U��)���͙n53�b#���'�B�?�T��lzi���5�턊:�~��y�N>l)����?�1q_! A��I�@��5F*��.]����g�*�E��	�S� �M��NS�ܛ��T�7;�A���gs��G��+����r1��)ꌵo	+��ba����;�N�CA�=�Nu.�oo�լ�Ϝn�$�r&��r!o͝���Ȏrҡ&y�]T(�/d���cb�8�w[����"��	��G��_�����8$D��zD�ͼ>%F����r��I��d�u�gҘ�[��߭ ���O�y�k<�2��냟ĵ���yIUk�t����z�̫�|$��L$$}/�<h]� ��Џ>q'�~f���2[��o��S8��Vڂz�w!MIrl�]�D�o{�=�\O�ʊ+"h�t�V���8�ҎXGs~C�BQ�E����{����:CJ�:Zv����VдP���L����ջ���񉈸��2�s��>9�`���W4�m1���C!��3 ��8u��b�o�h>ͤ�#��*�6�A�Rc;��Hz�����0���^�ۅ3�.|�}��U��@��k�z��~�Ŵ��פ���{�Om��Q1"!Z�U��l��y���*j;�	s����f?ᷧ�g�����0Zok1D��r.I�����ܱ<T����&���\_��
7�tj�����H�ڛY�����M�!�obzZD\�DI����g9���?� mV2GX�աx�vmӸ��$B��^t1+��EIk>|T�S�}P�/�J�\݉�e��]O�	��g��9[��Z�d}%�����
�w�%F�f#��fC.�������_Ѳk�Ul���4��~��C�9�|�e�fb�UN�iT6�^��q�×܅� ��Np	���m�WI���;䃦K�^N��7�)�F�o��Bi��"��/{� '<(���N���1Ԕ�8q�?�5q�Io &|���T�� Fx��B��pME�{M���n":����c��%��_�T�����-�d�
G�� �Z�g��f`��"�r5�����V)��m�n����.to7iI���bH��l��M~�����AE�P�"�*�M�ҁ�|��"B�~�T$cC������d�����4[�7���҉��X��~XCj��a�h��ᭃA���xv��ӎ.o��+��ew��|��;�4��*˛�������y^)XlN�Y�^dm9��y{e�������}���@���&Wߏ�qŹ��l��A��T\�I���Ø��ـ����xZ_'��ʢa����|�T6��W&J�H����\���eX�1@��`x�_�*�t�2�21t��Q��h���ô���o�v���C�'΅_j:�5δ ������es������j@�Q�vd�y�u ��t�q.���o�A�h}ҴV&��h�3� ���""����5�0E�(N?�	@�H�|�>a1��M�J1���왥r9�s��j����Yc���Wˋ�3�.x��}�}��Y���j�ɝ��5J��$��%N$����8�;���S���b��
��"۲#u�9��cSV�ٴ��5��`^�Δ�|Q��ōǥ3i���
�3_�,��E�D� �1Q����x�T�{�sq�}$"D �x*����������c�ťZ�݇e����Y�w��_A2GG��]@�R�cn��~8ҵ�!e���M�e+�;܏�&�F5Ez����gDU���4ƅ�P؎�8 �[�gW�6h�c"k���(�����{�-�.�T�ŋ7	_�7	���v9���y@�|���^I���Ck��oZ\�q�D�o1n!d���W�^S鑢T�j�)�i��G�w��\*}�(b ^�|�×��n���=��k�2�
���M^-b�^�3"���"����`�G��<�J6�{К�HX;B\���[k�&���K�{�b�R��'v��-_FK�ѽB&����ۜ���c'Z��jԊ����jԊ��R TrUO�P��H�� �-�������oz/�,���c����T�p⯥\�vB̬4��'K�}Y5�����{Ave��;�i�Z"^�O����}�������Q���jnǽ
d?��To����z��򁟡���
\�-�����(�ַ���@��T|=751��[Z����,��A���Ȫ��ף|P��CŢ�o�\���^�Al�`�'#�[��ݲ��{y$���'�
ŵ�D��Y��E�O�'lW��+c�Ǔ��o�;)�R�Ë�z�5CC�M�Ê��8-ҵq��Y`��d�b}�N��)`��j&�b0�?#��	y�բ���8o7f�ߚ��̦��$��i�����L�3��*'u��o:�d��2�Sv����u,x\Y�l�h��ڸ�z����Yi�����(�6��]���W+p���)t���x�s��ܛn�n��w����Y�g��Xe)�fJ�z�=J�=\��D��/0_��T������㝯��@A�6k��^n��ۨz������I�l� ���ߛ����� ��B��䷶g����0���NoT�P�B<���:�1~VЭ��ԼÐ4n�!u#��S"V��:�k3^��Ǣ��Ƣ����]��ޡK��R�p������h�-��nG�����]�#J'���*�X��,���~=
����q����Z��xk����y��O"{�z�8g=m5l�Y�R�0�B{�ڂJ���3ni{��k���������z]�o�(���-�ԥ��r���&�nʫ�{��]�fJ���R�0�~�^�������)��M$����&�R�
�8lhs��)�l���+R0/�Y��������7cӑ��z�/���mIY��������&#����>R�O���

�Es��	ͤ��Q���r~ژ����X��S�M�lF}�� 1��]�n���!�� ��1/|�r^���[��� ú�6_h��T���v*�C'?�_����9T쟹���؟\O�����
� �J��
j=V�q�JU?�V-7.Q�BJ{7ud.��m(��l���Z��O/z���6��5�jc���I!�"AL��]�s�s���Jk�"�w��	7H?��ysqY�5Gh�;�[��H�[�6P�2kq�H��{�u:��_�1�آ�:�u��y�3��1�h>k�?U4} �A�h,A���l�3�?�A����'{�'���n�̏�z�ʗ;��F?�z8�`-�ש����u)Q����!f)?r���G2�)���b�$bڀE�K���vl3H؞�$E�y���Ǘ�EF�2�;�^S�/�Wjض,�i�!��N�rVMʺ��+��<��� ����mRHyѠ��YY��p�u��a~�,�њ6�U�>��9��ݼ���-}��h�O��k��M��?�ve�ܼ�! `e�\�:�)W�~�8��I���zǂg�KKVᩦ;����賲2��[�V��ط��	[jLM3����0�a%٢ϭ�JT���X�{��%�����
��ϯBh�n�rAj�S�==!�<����!�Vġ�b�#�;��<���6���R�3���"���F��f��н��wc��jGdXiT\[J��7�?��90����ɑfptS��U�$����\n�s��<(IH	�F8C�O<]QQ`ePG-���t�����?�n�9�e��s�F&���a�'����/l�:~}��bm�	�~�����^�muc��L�� z��#����|5�vy�"�X���w�V���< ���jD��	u �W#���龁j��3��)>?�W��լ,{���^XKx�<�*�^�zC�	x�n��ʮ�4*|�j��]�y�h�*��41Ū��`����ث�#�vȺg��d�)����~W�3��i�B���^<mZQyҬRѿ�2
���b���Ք����a�}ބE�����K�V;��bi� #�=�HX�-94���3L��o/>^C��j��_��Sc��Pͽח��5W���kio*��F��ҕ<����A���E���R�	�í:�tZN?�-���QNh�0ߺzc�t�a��a�'{�V�D ���Ƨ~�?�_��}v:ͳ/��x�l����9 � H���g�%��]_{t�B\�}�jKL~	��-���S���DAi7�=J�q��4�L��1n�+N("�b!���AN��u�e]Y_K����R#&�hx3\) �,�Q �[qT~��_�/��	�{�s�������-r�dn�5@��I�b4��������L�E����R�g�~�Vo���� {tP5���%$�����^�+����{0ݫ�G߬�i����$	�~7��
�E��Iy��d�07������Lw��A_e�}���/kub�������1���̝呀-=v1^`������������X|51���j��}z�U�7P���1ߧ�!��*����P��첤�Iv ?�� GH�;,�,	
R!�0�~\�ꎠz� )��n�;�_W|
����N[f.��M�;���%sN���;�9ժ"6�ǿ�N�f�i[Ym��v�,�=Bwb�'|(ܟ���tU�(�t�|L�������-��+����⡺�{\��$�3a��}����1�V����g��r^�������f��^t��"�c��#���3�h6I+)���ɑ���	J��f��O�+r��c�8z�t��B�kdY_R�6#�}����8�P��fN����X�S+���[�݃ʯo7ˮa˽Dl��0�g�ʘ9�;v2~�#]]�o���q��ܲ�n��SJ� �u1P�Ts����w,4y��G�|��q�E�(�	��A�,�������M��
;�̤,J�ԁ�'��dHO�x��U���/vޚ���:H0�����G�M�a�l���� �)�8	j�s��-I�-�.%��ߓ �8�1�&���O91�m	*S��s4L���j�I�s}IAv��^鴷b%�_@A��Ϣx���2����W����z4�d�j���T��+����O�@/�M�⣚�����B{��D|�"��S��d���a|� �;d�k@�ߪRux%w�ޣ$���5_��<��-8�����_^�kzt��i+���>�]$߸�sv���Q���d���{�汳h���LF�?J� �������
}ҙ[��b���"&�:7g�O �fp�Б���]��c_��5��q$`�0/!�A��=�S ��% KO�^�VE9~(�#��	oҏ8�˞�sI�C;��v5�y���x�I6��y�*P�{��Cn�@X��J������쏠>��g*�س�/~��a@�ó���*�'��L���b�g>�>y�j�>�^x[��z�Y�,��թ��[�6����Ԍ��m y>���4O�ǕZ���� U�������Y����F�1���6�Q��͆�)�ɗ��~H��'��f=Ǆ�ӿ_x�����p�$�z�eL��2fן��ٸ�J/@X�
Bx?$��N��g���!�}���i�M)t8U�(��^��Ͼ�㯴��|
vT^r��!�������۝/����>�������������IK��Tq6C������C�^���?h��=��3uchQ�rS�~�U��~��K�3�ۮ�L��X)���VIZ�"���C��☿�x��@��-�� ��7?Ջ��Z�\��}1��U�9�I��V�d��n��4��HD�	Ћ�p�Kzs}��i���aXd?��\D�j/�U�;�5q�mSg�����_Pi!TB{���_�@��{#F��V^��� �c0P_vc��^ea�lWȣ��W�;�z�Jb��7j�� ��_�f�ׯ�#�n�	�8�ǐ����p�]٣�j�(��Eٝ�|�4��8Kr�����S��eJ@�&p呿BթMVK���m�������~H�oU�ھcz�~�	�'3Ё�f��!
�d�sb�X����
픈)�L�aw	�DMϰ�a�A�<8�2�k��"�ws�F�du�����;����E%���O�i���_(�=Ԝ.>��|�c+Y ��E��R�k}a ���PB>�|��
���bR��P�z�)?9g;1���r�H����
��܂������ݙ����A·a�n���ֺ0�Ĕ!�GL��(KcςA�S�ȩňR\�yY�_��G��8#��9��i�ӕ�����G���	�ƪ���t��sm��A@���S�+.�	R�FƻDך]��z �E��2�8ҩ��Z��B�_Х��H����@�Γ*D���&r)R�{����T�_�cV�Y��T��q-(��� ��DzP�I��t)���k���B�t,)�jP:������~>���7w�̜�+sgg���ma�i �Tk�ɮ�����аu��9`lo��/�9n�{�\%ċ̩�L��;W�6h�P{��&��,+�PN�!���ɽ2��͝�����S���Ņ_o6�W>�^��ڮ�Rқmp"����_���걺(s{����%μ�=Ӆ�k�'�oP�����Uh<�m��mi��D���6b�J��Ȇ��,\�	����	��X%���W�l1�y3n�a6\u/t
���nx_j>-�2E�����=�*FuM{�lS��j�0z�|x�	�(���Ő�nGe%eph��}]v��w����&�}���oK�X� ��:��܁e��(����ZAT���
+��� }9צAT���;�An��G�x����7|u��
�g�E���]!��9�}u�	M����ɬo���~����'��E�����z��#�n������6G��^ͳ�� 䋇�0�q`x�w�b�!���dV�����CŨ�kk��Z�*2���G=�ש�]����;LVd:J>z���x!ס�%q���3���)/R<�"���(]JI��f��o�Ny�1��~�ވ���B������������v�~h.���AT��Fr ���2Vx�Щ!bIK��<�Z~�刧@����C>t'C.P1�9��tsfY^�ѥQw_������'��Q��zD��~���~#�I��/}�kO�d���j�=d`�(�bn�ˎ��!��~���9t��M�)o�0@'���l�sq�j1��@D7ᒥ��Ѻ����5� ��niOirӹt�*���fcrz�gr�5x;bU������;t�z��ջ�e^�Xf �#sH�|w�qxL��0�O|6 8U����C��8K <�7�8��p�d�$�d�<0��{+6F�:PZ��b��s*;�A���"uș�h`��(vV��'����e���$q �	�?iY���l���F�>����ymΡtb7s���j՛5�Rʡ!J�y (��@ݣ�p"Bi���A��J��g������-��MW���'�\�� �N�M�vm]qBa?���EZ����$0�JHPF#s�Y�<)4��ǁ&�ӓ�Q��e�ա��˶%b�Ċ|?��h)���7sC��㕂�X"��g��w)���t��i

�i���)r�1��x*&����X�I��<Jw��Z	�U�;R������>Q�=Ӂ�h�¬��*j���c�y�+}�}0'��\�H��e�t�ic!�¬��R3��p]I :i���zms��z�&�K�g���j�z�J���Z͝��UW���19<$�ɯ���a��,�hiqgj���
��(��s��Q�&b;R�N4p�,������_}8\:=�yI�ۜ�P m>�\�9��&(���]���7c(i�MAF>��t��?L�x�ut$�ji�1��鼔ה���%AN[sP��a2��?11�	R4I���-N%��ڥ]���*�˿�Ū����pһ�t�D��Ǘ�!ǉ�㴔����*y�����l�i��{���D<� :g�4�MM������5�oo���ݨ�΄��d�b��F�����|�+u6��fq��w��'�a�����6%��!$m��(���	K�X^٨�	 �������c�n-�����y�IfsOk�GI�g�ʮ�O"�9�4�����\� �H��f�N���H(h�	g6�ʹh�/��c�mG�U���a�⑛�mYG&/E7OOfQQ��]�:B����'S��'�]�o3	��Р�������6���d���g��D���~#o�ת�J�L�΄��6��A��4�$س,!-Jb_N��jl�@3�5�A^�S1\Z��Bx���>�u�"�z��G]�9�����[�8��hC��f�01�U�֦1 �3�C W�̉�N.Q��kR�^�&�o��1�6�#X		�4�-�v)p��ϭ"^���d�.�Tc��W8"�h�ۏ�6�2�۬{�%xmH��H��GGz/'��4�c�*4�T7.'e.ѿRmivM�1�k8��{q�n;?���9/z.�l�Ɠ��m'�]�[�EHA�եo� f��(�jN���V ���o���(`z�{߮/���4訕��>C�;�i2�i��K�Cݸ�s�������Sn���{]�ƍ匛��=M��R��bs�����cz��U�%t��Q�r�܊I���o�z���'��.���VJ wvԽ���=���J&�ӎ�܄�(���0�@�1XͅA�К���Q�R�&A��Άu��G;�K�2i����)S������7e��%)7��6�<���i�Pzy���,e�'cz�Ub�!�k>+�3M�1��j;Q���Zsw�=*<�y�R�o�jv~{4�4JWO5��Fr䬤�ZV���y+�"����fB1y��G�W�eגk	j�%Eh�}�Z8W�u�]��XB#rq���J���1r[?�:��6�m)|X���s�/�O�����M-���7��Ӻ��n?���pIW��3ߚd�o;��	�d$x��w�*�Rj�_J�~-�ZY��*�vݛ��j�k.��ʲ:��L�YΉ˥@^ƴM���S˝�Cm��B���0�����M`fPU�@D��I�d������i��2��Qĭ#3x��CD>"
�����p���gr�s-���EI���z��}[��s��4l�<�5���#�u��Zl����<�q)��`���GV�C5���N(���|7��S8�I���Ƀڛ`�Ԯ��T�]��I? ʇ�i��r�5e�넺��J��LT�����B� 7�S���=��.�]���ϕ(gc����.�e;�D�*�m0~x]��5�>.�nk��aa�?%>!�ډ�������]Q��'_w3��k��C^6�Y\ Uf��y���ϑ~�d�6��z���*#��M�u9E�^��[��ѷm�0Hc��n]P	�⭪�4��h_�dcb��{�НնFGU��a�}0��:����Fs}1~`��-��/�S�|��� ���� ��=3塺;jȣ��mpH��і{v�\���;�Y\���c��߃e'!w�w-k�5�nѰϏ<�
 O�{A]p���j3ָ�hZ��^�u�V�eI�f�̛��R}E���Bk�Û*�,���\�/PD����F���#}`j�����	Z�"�G�an3��
�'�r`������sU.[�t�!!(9c�铯]�����fb"��l<�~֏�4#����೵2~�mg�ok�K����/��ds���gq�^�M��窊�.`���{��	�k��O�绑�D'v��ߗ3����7j"J��0�K}\{/:Ӌ���ۄ��n;�����|��zx�C�T����.�A&���KO7(���_�wJ�=I}Z3*T��h�����,�ssb����R?��cG��?%U�L� ,,
�"{zT�(����.��`b���|l�A7��q}(��4��ͻA}�ќ|%nXra.B�v�ikC�,�lӊ�j��ى�\���kԵf��}��]�J+��k~A�+�U5eG��Y��mPam1i�<=��­����G)+0������+:A����R��m��3E>��zP*�����U<��w�5�~dg �nz�:BF�S�ݿ����,]=�?���Gv<a�oC)��%9���ujC#D��8�dʹ	� ��{ ƥ=���a$i\{���^;�x%�0n{����G���Z����K�4`7P��{?�,�� /��z�5�b4)۹)��{U��f�A���{>��G;��f�3l��B���E n?FT�Y��Y�p��*�6�6*T *�tmw�X=���x��ʋ~g���C3G�����.�q�lK�X�շ���xKo=6ْ�Y��2_���Φ�E��d��k,|xb���+��H�튚��N)��{t%Iq��_9�J&��Q�������{1�R�����D�@ݲ��6�7s�Ŗ�o�����-���)����7�Y��%_��B��x!W��F^..4���ř�z#�*�r��b��äT{�͜i��˩���I=��^I��R����+�����&t��[���wv6ˏ�8	#u����L(n��o���x��^�}O�E,���W]�~�@,���>��TPr�3�a�Cf�CtRThg�t����1���LĢw�O?`��ۣvY�� (-/�h��;&��P�ٮ}��� gW׬/?�-��۞F·���6�~�������[.�ud��'�؈p�4,��W,0rm|Mo��R�8��_���9�
�|�N���SM� N)T-o!i!U�Wv�*��]`�c�l4�ic��+y&�S�J��6�TD��7�^��OMSj����O�S� *�H2dcW�7��DHy����eI�G�1?�����t������?��)��1}U��e���{pL⛝W+�z�Z���5������t/@v�[�[�=FK�[3�%Ue�:vg^D��F�#G�ILl�k��E,W�/\ka'}+���_�{�)�L��<��KW��m~�!p��kʓ��5��Fj��}g(��.����P%���n$��̊�O5���ോ�?�z��	��O5K������L}zF�ݯm/�H��G��l�:ǥ���- �y7�u{�l��ko����p�Y�?9�o�s�W��n\�TYqQ:�y��A�y���!�,j5�ٵX�'h7����������]X�
�^Dqֱ�^�VLVH��H/c�sn�5��'�1Tޠ�lw��H��TI���b�̲*��R����._�)��AJ轥Zˈ�ZЙ��:���K7\V}5嘖���+}=Vq%�Xh}:�b{����w�'bb�_�mo��+d`Ž���6%o�F�m�V)[�fkO@:��<�&�3;��֒��c;�M��DzB�a�07:�`�N�.�Ҽ�����.ٝ�+�"#��d�ەںe�����R8ѱ,ꦓr^x폫�xz�"[O��Ӈ�y��&X��' �)�"q]+E��SM�q!k��f����)�]�Jc��¿�v���K����6�̾���(.��;.��ly/p{/�w�d���y'R�-l�b��|C/{:���u���^a���}�?p���J1����F��˧�v��:P5z���"wى�%�F�	�� �YА��ʽb����q����W���+�X?�|t�� �ڂ%F�H.FF���[��]�BU��/�M��������o��������hM�n�&l4�Aj'��HY���;���2{V��V�7o��(z�je�5�1�M)i0X ۸�I	�W�#�R�_r"�����F뮷Q���3�U�7��j�-/	��Ayej?�������d��I��P@@�W�'42�0y#��J�{Fq����w�[oa}�
Hk��>4F�+.�b�v�	*�v�f>)��b��*�sSUt�z�ʪ�*��b� @����	f�ZSp�^֧��]Yq�����N
y�F%>�[�� ΢��kØ�Q��b��IEv��Q;/�d�!/b<+�zk�	�
�[�ڑȠ�Qi~h���o��=f�D�Ӟa,�Bx?���e�7��v9ᙴ]Fd�<(��o��8�}�EA�|��ݫ��>抦��N�c�6��AM�v�q�cT�J�=�rU��z�v��^BQ��h�Ni�{lf���?~~e�`#�Ԧv;�WIv� �=�BΕK&�t�<Su����4<�Z���䡅JfC���O����}{��/����u�5�E��0�}Y���wjV��,.�|n4���g�,�e�=��)Ƒ��d���ȃY84k��0��#�A���.��Tg٣�(����s`_����$�\ ʾ��j�>^�/���+y����es輿�zЯ3,+�J;����QVw�@�:�C����nB��X�W���|d&*��9����mE	�p"?�P7.f]3Q�t
ۙ��-�vb�&W�;�����ixL���[�1~s"e{�����{�Ew��w3��
vt|6�˨SL*���>A��З�� �l Ԧ>�q��7"_��.�,�O#<,M�N�?ag�Fj�]�Q���ݣ��c�3Rޔ���>��I��饼WW��� ؅%���Z�t����/��(�4�Ķ{�c����S=}z#�Ǩ�"�A�`��8��tޚ������\N=p����]z:�Z9����x�Wc�V>LeNc������P+7����T��ڱ9�`�s�f1����H�jlQIV� ����>�g����Eg�j�CAX���\J�,�#�1�vЗ�,�ߵ]�,�<4���ݜ`?��gLl�"9�}t�A�e-Mu|h�UL�'�ϰIR�����K����i��b?Ǧ� 7�U��=�HP�������"2ϗ.;ӟb��� =�R�r	��<]��c(J�n6��Z�=��X�U�[���9|�7Z��x����ɾ����*��}���r/c��ն3�<$o�IO�Ib''�<�O�˽6�H}�H��$���%]�=0�T�9��� #���_����m��	��o���K��E�]�`p �0���a��Ny��#vQ�����Q���#�}ɛ�f�0g�赫����R��s�&<�]�k��'6t=`T��WJ+��9��I���_F��^�����|AuJ-�W��Z�ع����fB��JX?�����]x�A���Q�~.�e��5[Y5��QQ5�����y��õ �d\B>RX�"X��,��/����9�O�Ur�*�$_�)���x��֫���j�#���yu�rT�t���w�3��BmhҊΩh�%B4G��8q:�8e|U:�K1�oN?�X4G	V.XbV,�o��;�č�q�ot���W㪈u��#�JT�z��ި��8"�{G���j�Y�?�~�Vw�S��*�mOKUy6u��F�<(-}���j���0�R���Pc;��ٌ�}pήg8��K��r�'�Б��D���h9�ta��)-*-s:'*�5~U9F6���d՗�P1Puxs����o�/�H(f�������ր������< ��e��<���sA�PxR���=)��Y	�f#X�U����6����BK�[bA��+���M�.���}d=����hNd~8�軆v�|��V����e�J&�4���". x>�1�
H�"�P��!������]˗��t���w���;��Q�Xw\����7]�[o�ɤ���B���4��MN�Sw�΅��i�u���彧Z�E&���U��	L����n��G;-�f�WQN����; Nj�E�P?���{��?�ON?D�-b/�<K��ɟ֡��8R�gC�����a��y�׋��8!����vo���z��,�
�R�}P酻k��s����~F��]�۪H(���n� E��>�S!�8�h^ *(��v?	r��&�M�K���H ���V6�b	
ք|��������N9���d*�wCg^�v"�6G�kN�0�5�F|��&6y�w[����&V7;�c�:r�*e[���h���F�_��mM��=��cW��$�����W��R�~Ȱ�3?h�������k���I��<M���Q!!�2�k)R�i��������Vp�j��=��WRL	�zX�لT ]�m�Z��LyM��J��Z�Eɂ�~~(R�o��)(0n�v�9��77yU�G�>3�]� �Zj�ػu�U�8�����iP���G;G��r����&�MefM�N<e��SM�u��]>t�����;6y��bDo\ �R���bc%�b��+���>|�k�76(7�����]��W���hs*��.�q0008z��I_����e9�,��-��9i�37��m.� �@�'���0�m�MS�er�ԕ+/a�������N_����/��
l�kœQ3I�^���Rv��d?t���x*�oi���w�ҝ;U�;����5�.����^O�u9+�%|���T�fd)��7�7�[�i�J���$`���y����x�Mwж�hX0�Q�Jp��x��4��Ɛv=��d��6��ݍN��c�~3Q�dz0';m��l�W!��aO��\��*��a�ȗ��$�_p~�,�Ǫ�q�*�����p�ϕ�Z���'����*���ZuoN�iܾ7h�gr��=�^9դ�ʼ`3>Y�"�R������{���c-��qoDġ��L�n~ؔx��@��j�d�����zm;�j2�݌vd��Z�"���9����ߨw�ef��ȼr+h�W�b��+�n���MH�F��\h[�O��;
_�`�(6����~�n�t�B�P�4�<˚s@~�cC�;"���cX@�ռ�'�P�C��clh���Fg���5��ψ�f(���/�9��G�q}��K/�C�kR����=�͞:ޒB�%�-�aƔ�tM% 4��D�_7�x^*�Y��K�ڧU�q��?�`03�o�8?z��Im�w�Df�ƭ!��QA��浶>7��1�i��5#+vl��Sor
?(��<(����S�z�2��5�#��B^���,���V,�~�N�~�u�,y��;��TV��Z۪��P�;�u��f��޽���1�h�F@a1{�l��[d�-g��? U��;���n=w�rk:V;�����7>�uS"0,ƨ�a;O'>guz����Z���O�j6|\�m�\�:����oAv�������+ZH����3��-T%��8�׵Tލ1�n���Mx<�0��j��/N`u�z�*_V�ap*	���)���4��;��`<{��+��o�R��g�}�7�6(K��ě��;;�+	Ǉ5�tKC�E�7J�#!�Ү�b�i��Vʱ�|�Œ�RE��QOL�K`��ڷ���$:� �}�\thR���S�c�n��)#�?�芵��h5]�g�\sv�!KsX_��Q�L�K��'�u�z
.ٶ�zA��D�|�����#ѡ$t��k�I����8DF-!h+��|�B	kk�G����|^é��]o�[���V=�|���\J3� u�}sn������@!;��lш�z��7?$�3�A�_�rC��qB,+c��}7j�Y�{���|ӳ%�U݌��#�>��K|���B�H{��變��E;�[�h���Y��:H @呓�gt�=$�\��c�DOx�P�����R"���t�o��|U�EWn�t�%ߟM��<#yfiV����[����^[���ZKY~n��<�t���^<�3�Zݹ��n7�θ�MU�|�G̹(�{{4mk^�ڮ����9CT�`lmeO�����=s��0`n�<�ߥz�.~�E�O��뵔?�c��q{�)��$�y_��ȅQ�5�8얘��]� <"���>?I{6�(k}�hPS�̣/�$�����jrZK�d��-'��1�š��`�9U�U��;�+�'�ۆ�X��Ee�<a�ɏ!�*4ZT�9i}J�d��G#�.��-s�a���h\wIP�O[�(�O��**�Ox�]Pʾ�RZ���{��k�dO��>��6s�^^�Y[�;�ކ6�"�I��33\�k�(�jϬ�׵��%��)�ԯɩ��9"���_�e2:&�N�K�>���P{k`J��	��e��[�U#�{�<S��������c���L�'�1�`��߅TeVVֈv������O}3�9��i��ݦ�zźN��]�\zQ�[�ԑ
����2�p��K�����m��>��#����Ǽ��p�y��i�P��̜�y���9������[�7�S%�o��|��nl�O�=1�rX��jﬥs�dN���B�
�@p��v���\��1��se�$��-,<� 1N�qs�{߈x��/��Qa$irDkߩ�m�o���y�ɰR�M�Gilě�b�k��D�Q����;N�.�n�uQ���I�\��=�3��be�����3݉UǶF�����59Sϯ�;3�Z�y�����}�q�o)����<HH��w(Z��O6������q�cf��}O6
MVHd-e ��5r������\�p�y��yGt=J=�k�v�.B��!>d�<Ē��|�#�`ͶLĆ�u�[o�V0�s�����=�A�F]��̹T������],�C�����=��P���N5�:�y�g�[G�QR%&6l�Mݫ)�Yr�z_A0�Yw/xՈ�Y;��e���f���4�<�e���p<�'9eW��E�m���\���͝�HI�1�)Q�!>��g�]09���|���kw}-^�-���vZ�Se���� )����B��ٯ�F�^E7ښ!D�W/bi�����q3���$���b����.���Qʆ�w�5�}hZ��VͿ���pmx�����;��J�����6=��n6��m �Г�d��o����I\0��%�[ڦb :s���+������|J�hj���%h�Y�O��:�����ߊx����=�Z��+�x��O�o����g��5��u���渲`5'�%����I�)���Kځ�-
��LGo��	^�Si�~a�3�^AzZD���Þ�"�&��wN��[�>�E�'x���]�Y=��"�!۬�J�_�L��15X�;�[y�B~���P�~�D��;wT�S�*���H��1��T�1\*S����t�L�vvmj���+(OD[�o9��U�z��i]Y�2��9h�V`mN�奒��k��ȧ�{*}P��4jh�`�����Z���D�pQ�s"�ć��.�n:�n&a��V���435�<�(������i9�� /��yD�l�j
"-�CfZ�o^�ߜر�j���p����o|c����{�.Ъ����։�y�&���1���r���7Cf��g��Ĝ��dK���̴]AU�6��kvW�?�'���фv- $wB%�.��J�����!u�7�~�� �Oi��L,�9'@"�˝�H7�����/]N}�6a��?�*�j���i~fiQ�Ҭ��kD�8/����&̹�Zp�� P�y�|�8q�p�̒i��o~����.��1�q�$�T�_����>�òk��l�v�R�W>�ab�CT���Z/i�� EH�h�Y��*DQXH�0O�$��=����.��;��/M��kW�׍l$��S�\H�`��I�, �0Î�+��.s���1�v�b��{�]|�ͺ_�x�-��GE��d��+��*e���U�Mk���������9�+�&F9ʮ(Ä���yy�<���?x�q�E�^o�n=��}�Dۺ���n"-)�'���\4(5���%��,l�˰�~�ڷn�p���u��^�p�Wો.�@6�����9��Q��ӊ�PfZ�i)WL�2Ϲ﵏k�{�����-Z����`�L�*FGB��uz���uu��nhe-�S�;H�\O���N�]k��r�o`8J�,O�����K��
z���h�,������4+�x"���W���Y�>O˹*|��G��[���b�J�Y��ɇY��w����j	�ܪ%.	�\�|��1�rU=[��!.��L�n�V�'O�U~F����1� z�Lohol��4m�ݔ<���ѡ���KA9���h�h��nn�3��Gl���H�"�� 6��� ��B	<���h�4�Ý��7�&�UN=J�T=="���;y\����:.�ٝ�
z��<���p���4s�p�n�}$F�KZ��{4uA��U����]�ڼ�&�ؤ��Bp��q^�`I>9����?1��
�+�sFK��Aӏ�~�iP1(��a\�;�{�?�0��O�'����y����Cz�x¶��%�礀4C�Wh0��^ J�E=2�y�#�垅f$:�=*C�o��o���F���:��u�TT]�М��ǹ�/#�*)��k�-�/� �Xr�D��p���Eo��Y�<����?B��Ñ��������:���R촀^�i��;�j2\�	Sh���HN�uKD|��+��^QQ�'�'��<c��Ăw}��	���2�]�ӄ�h���T�F����
[���S�=�_���U.j��H�&�?�g?�(��]�*S�=�������ζ_J޼.S�c�*u����Xc�TTRA�����^=�����$E!�
���{(\�f��=n8�o�F�����&�ȶy̛q�����6q��O/(*6�Y�:������̫qlR�Wz�x�qyV��p��I�Ľ
��A�t���#TV'�3I�_C���U�,wÀƍ J���o|�0��lK�D']S��̦�YVe�Š���7�/�ʴ�)-�C/�陸Su����md�>���>0�l��O;C�
�Z	�QG7_�@��Vj�'�Dce��I˨��M�rQ2��c���qO~���^��J��(���3�TT��pLq���^����n=��;��h h�mQP�K�	�Ax=��6���G>|�I�3���Ɣ���^�S�F�<���46�G���|�%�o]�s���3 
��| �Lr��L�-z��>&����_B�ۗ�  C��ک��Ϊ�0��EL�)�.���Ɉ-.C�-�i�@F':����ƨ�$� � ��J���ZV/�\Գ���_����s�2��ˏ�p̍�8���+p�����а��X�m9_�%�o\|<���Avv6?/o��G�3}]:�������+h���u-廴�]��{�������rtKV��c��7nD̺{a7�]D���,,���Bm��g�3��v6�i�ж�e1BREE\����{C�n����yy'�3��C"�����6��
	i���989�K�ZX�H�����"���m�h��B^��y�RMEE�߿NOO��a0+'羒����{0x���W�~��&��B���J��aHxv�!��i�"���v�%�4hgoR���	�w�u�l�%�/1-p�Gy���u�o��P���d�>׾1�a�^�����N�My����:RdV��Ξ�JG����_:����.��Ǜ�3
в���L�@�q;��U�Ik��ư+d����� ��B���WĞt_����6�h��I2��yOy~�7۴޿�;i�s~�3���u��]�	U���9k������;S]��g�~r�L�������Zn��<3���5=����v��Y��"�6�=�JLY}z��sc�����S,7��egn?3��Ԓ'{^
��/0&p�o���8����9gPFE�skm��LJ��Ȉ������Gk����wWrRд\e�a�>^Ȃ�G��t�x�I�`;�s֔\ԑ����c��TW������}�9���З��^;���f��}'b-f���<X��-��x�ga#+kxo%!I�9�֭[�`	��W��|{}e�!�����q�֏`cOmuuLv�%|�K�P�e1��HVI-�*����=o �o������Y3�U+��=@4��$����8JA�0�*�+�����2�A�S<�se���/����9|�������_���%V���"_=n8���Y�l�]�V����h^���I�yH���IMM�f���fE�����g3�9z��$��_��uH�.��A�:���b�w�DӪOQ�Q��}�r�ܧR���sb=�d��S�,N�,��&ưȩ4�40�ȝ�������=2i�0X&S�e�Z���D=�������G/�����n͗�����,��n��Ó�  ��|��)�[��x.*�7�~�b��%P��#F��`�⛚��w��������a��	���FEٕoא+mS^2�D���"Bq�V�핐��X��e}!��Ut���,t��6#�o"���~0v��$�]r[��^:��٪�~�U�);�՛�u�"����rW�,�zՅ�q-n ��5NQ���q�f)�LN>�]����
��|��!k�-��x�툵���Ǵƨ�*:,�Ý5[��.�͗B�ġ�w#.�MÕPCg��NS�����,�uQ�7��������� �4;����޵��h03^ �F���ڷ3FF�s�v�=1���i�S=�J�I3I���MY4`��"���u����~���d�F<���U ����p�1��))$0�jƖ���B���l�"e���#�}�ݗ���/�e��`�C?<n��>�l>�'&�=�����V��8�&��/ls��N���ަ�#bb��IH���R�o}>����:����~�����hJ�=)&`�_=�2�Of�v\V�����%� H=�l�8�*���<!�#&�^�X��<Z}@����K~u�\`r|kJVJ:S3O�zq���V���30T�Y ����gsF\�l;�e�
U_�������Sj�^�E4���ʯ�Į@������3�n�е��-s�1B�Q�D�N�������=Yʒ���Tq�Esy����uY_O4Gbjf�
�k�F�I���jA>T�H�*B9F˱w((脠e݃%�f��R���m��]��5��9d��g��0@xE�(�*��a���Q̟�݋��2_�j�{��q�e���A��_^�O�@����f� n���L-�ߺ��͍������������B�g^�Fb�n��V���\�P���]���I"�T�BD�-���ݕvA���}c{��>�	z��!w�䓯AtC�H�.J[��e#'c�/01�كygR�Ӯk�|�H�m$r@D-�MM��ӳEU�^�()�@S���;���L�؇d���
��%k�Q@��i�n��:�����#���ϔ����b��� Ҩj�]��������!@��ghɱ�j5dy
�?(�'9�_&T��H\_׊ʼ��9� �����Iu�,:uޞ��K~�\?G�gw{U3nx_�Hر'�����7�  �ND�L.��X� @W_�%����Q��$b|Q�p}����ݒ�u�P�/_?���/�t����qQ���ٜ��S9�� ��뾅��@&����O����S)�E�q�x7?P�<�CAӉ�h��ۤ$�mUUU����!�6	����׷V�a����'\^��fw�_3dH�����,f:)[cf_1Y�T�J�y��=5�ϝ���x,P����;�q��-A�v���OiZ(�}m(\���RݪV�����7������ogw>���/�4�4\�z0n��� ���4P�Zh�R]迂r1$9�<Fuf%w&o73�2�a||O��V�,m��ddmk|Pن�V�} �G��� ���(:I\]\\�����3���� $7h�z�b�'+�9w]�秣�o�� ��e_x>W�Nb ~�$bd�N�ɟ؞J  \Mc��b$t�6\�8��n���\� �)@k�'ZN ����V��E��e�b�\��
���!!Uv��+m���l��Q�@���;��6��2�����7
��.>kpf2L��%��:��U��~�J R)�)\5��������?*~8��DFcs����'�Τ��}q⸴�d�t��V�=��M�L�V��r����n�� �rp�--��v�2�h.��u��r[ �*ㆣ}��Y䍩��}/���Co){N��R�R���/��g����~gV!셥|�z.�T��=>��Q@�z�B PD��up������9G���1��#���K�r��H�o��қE�%en��M(@ͱ�*m�%���l�Ѝ�������k������d��ͬ΂U�z���K�+���OSM-LKv݀����R'�ƴ79�^n��6�uA�[̯�T?,�<c~���C[�x�+��X���V�NG!�tI]q]��1V�E�w)���,)� �\����m�Sss^����4'�ϓ�s/���R����H&�5���9�s�{PP�T��`�+�'��ʔFR���| �YݱSj�tr/��;'/��=R~£�e�*] �U���w!us�5�)QG���������RO�8��Y�e�>^1��6!��5s��LZgh�F�^��tU�����;Δ3�M��]�|7;[i�1�p������EL @sc���Z�'�	��~zѰ��>�LǊ�L7������f^��f*�s�+������&</��*O5�=X'7K��zv��_����X���1�ݱ�v&8�� 6�����b�i~m+Ȏ��	R�A��2pp��mB��d��݀�w��7�n���+2��5�K��h�L��zuoH  �� $.����@;�;Ha���G�2_6����駓�/���3q�;���n��������:���hbnm~�Mε~�6�f���'#;�����]�qqs��"�h�����=<Z)��(�w��Y����cae}Q����������J#��N-��8޽�,R���_��v��v Y3� �Cd��Bq2��ܯ�di"E�	�w-�+���|�/%��9{r0�u��� 2�]���3�}�<f[��'�5�0xئ��q]###��
�����* ��~a�0zqcK��cY�����<#��� ��]��dt���	O�x��������/p��Ї�B.�AԜ�:��]�CBkp������e.��̒���}������Į)����Z�i
�y�.y�B_&/(� �t�-��شr�a	
�+))]Ѡ��H����W�!R�"�<r4��}��*���ʝ�t�6+I_�p��V^���\[����ﳑ��Lw t:{��S=�޴��k� �nqqq�4�Fr fF�iY|@'K&˹���k���x$W�ƱRI8}X�'���-�+�@�ef����ƾVj=�bIE_�����Nof�����K
T��r۲?|��a���*?ڋ���Y�񯿟���&�{�ei�V�2
ǣ�ɖ癘(�I آJ$qP���]�����fŖ�ǭ�0�7~���S�����w�}&c��W�>��O�����c1β]q��zx�+�`����{�^m{ܾ)��~J�����:_B[24hK�4ճ�߽~	s�����S�P�I���%�����P�Bh���X��)?`x+�YK֗F�響�ܔ�<��m��`���I_Da�u�0��	@u&��䁍@?Q9=Z��Pu��dy��������"�O�h	5$��I&Hnj��t��鿸�,P7%�1�Yq%TT���?��+����nX���g�±�e䌯3�����'��l��+g�-�%9�]�ï' �X3:ݩ+0}ţ���Dq�Y�R��#6���Z�t@~�iu�.R�Yo��cc�
b��AH*���" �t��t,�t���4��,�)�  �,����������<�^�#�}��9s��:�̬{��9!C��Kh�^�5�~���t�iy�%El$����}���Ra��[	8������k�P���2PF�q�=P8aR�.d��SRQ�ȉ<�~�VX9r�^�MO~��(ͨJ;�~�OW��H�B�v*�� ���Vڊ��+��~ś��_{>@3��.QWP �3�D�L�5Ͽd���FR"|])���z��3g���a�I���$���lP�.�~�d'"���e�9�����>oߞ�9p��DF��S۟٪���[9�cވ�ϥoNd����3�&�$�7�'JX����KSc�%w�/��^  x�7r��rݶj1����RK��tvvv0�!
�
S`1P(7Xl�$/�g�öt���'��a:�}�yˣ�",�l�T;#�aa��9}��
�-��h�]�}��aG�B�J\�x&�ſ<������er���{�8��%�[��$���`�+����9�/,w'
�k9�`�����{OIG���?�^Z��t��yҙ�\Nm�e'S���E	��y?�6]�d�w�-��GQߦ \\&�؀�����L�䚪z�Ȝ}���Ib�T�3h 2 SK�S��u �eF�����M�^�h�����"9�'�$<�cSA�L�0��ߐ�[-�k�@v�$��Ԓ�4�]���'�4&�����m�T��E�Ԥ7;6u')�^t���c3��O}$з4���u�� �#uj�q#UP2 �[ZzzC�ut�������+TΜ9�^�^e�4@�NLz���cxfl��ы[���?g-!�vl��D�&���>�_��(ණ�a$L�>�Z=�r��
ݛ6_\����l	���oZ7R���7ByH�pEI�V2���
�eu��!H zP`�<Ľ��ςp�.%%�&X�*g�����J��['�/>(����G��i�d2����^�]� �\��,��0Չ��z���I�꒧��N��(*)�f��u
Nǩ`�����G�{�0��&|}?���ßZP�:qq��I�* ��h��f����kY�@uV	/��=n���MG�C��a������;���j�/ba@%0���H�T:B��3���"''�ܺ+F�) � `!�?���6���l�_߼�"۬�{s�ɈIn�y'v(W3z��ŋ@B���������W�.}_QML��3;F`t��K�Hev�o��Q�^�}��/�x�����+��`ھ����- �kX���b_d�	#�]����А��g�$�U ����}�"�ϡǢd8�T�ig�!,,*
�aY&b�V�\���+�t'�Bur�]m��ҷ	�}?��KV��6��LN�%4L}�C�ޟ�6|��Ý?���]t���w�`OX�ss;�i�nݺ�f�B�,��8@\M3�(������O3���p��J��ˮX����O�z�(/ �j1������wG�!O�~�+k������Fh���c���Z�*=0Xc�P_2=Pq�ߩ�@�I���f6�%s����a�4�!b&�e+�R����Ȍ�>UN.��(IIv����(�=(�S��k�&�� c �p�9����bD��0�MK	
�V�O�"�v���(WD�i��	ȷ΍��ͫ�|���k��P�����ǥÖ߿�w��mE�k����֕��+�W���+8mg~�ߝ�mWZ�A#��JZfן@�w�л¬�oM��a'�|4�hY<4|G��U�^�Q_L�5�7J�Rd�:k��v��N���S��OB,��^�qc�����2�|e��d�/���՘��J+4Y��-t�,�~F�9O�]�h�'����=��Ջ�j������壍K���&z��ΟD�gإ�bB���t�ߜ�%�+Ӝ�O��;[$�5�U���;:^��Hd���i��P�@_
�@+��:�#!)����ߞy�{c#����8�z�2�CtqJ_._`�uvb���1���J'�l����T��h��H�5��C������
*i1��G>�Ij)Ht���u��v��Q�BpZATS�y��2ޙ�f�%,��U>ni�d�S݅TB�������rZ�8��P�5��q�U(��'؏s��S4��P�\1xZ���5����0cw-�qz��~���fʀ�8k	�8�k��=eɟ޺��#i���2V�q\@O��S]��U���\!c���AHFxz��3?��΢!�U���b}��wg��~�Ў݅&��"3�-��f��nh*  ѡ!��\��]$P�SI�i���<�����8W�5�2�_�\�h��C��x������;�+y�sa)������R����+�,��l����[�J�A���U�H֒��Q��N���~T��;�-�V��G�{a11C)��^'���׬�&PO�KrM�q!Q�xp���������~ѱ�������|q탦����F�!�a�����'�3Ƹ��斖��x >�`�
M��+��$U4�Ed�}K�]�0Z(dAF�����c��e�O���6�N��g h,�7E�RX�]�Sɠ��kx�%V���K���ʵ����O:o��@V��/��C&�F�g���g�|�<�d����3�5��lv(�q�<�ۆ]���`��X���>s�,��uu�%�`�B��v�g�խ"R޿?��WJ�PY�[OO�\��N�]m�����{s��>ù�.%��1�����ұR9?~���������c����/x�YO}�Lfy��e����䯆y>���[Ho���&"�?�B!RqO�Ľ���f��H���ii�������>�O����r�>���v�n���I�s�rt��4�y�QO�=\Y	�y���N;������@h��Ŭ5����S�Ε��.�i?�^U�J�A��T���� ��۳)$)''��{��-��ˤ��|����2@�c%Vug���x0��#��Ā�q.Z(L�>;��xf�ʀ�Pcm0�a	=�PR�BT�A�@��b\H�8�����Q6$. ��ߔ8f��U�D�c
����Bw:��8�{+59Ef����C<��]�lnܱ�AG�w_�
E%��?����]ۭ����
]�O?��V��J:z�Fy��/Q6������H���<�X�\G"]<�>޵��5��� ���,�ʓ��8t��LB{���p�7_��u�2W�q-�T�Ş�x��ǵ�Bb�䀵f���938%=�Y"��pG���]#<=e�����7;�2>y�����²v�
n&]��*��\�, �����.�TV��+�!$ t��Q�����GyZ��r�lj§�~��~}�I�+��nЩsĪ���a!��S��P
����8&g��������U�a
��]��@K�ڃ��eEDDBz�b*�֙Ɇ�]��JB�;1V=Jg�p~�Tw;L!�Um�{�Nq1�R�c�8��ՙ`L�q֑́�wҸ��Y",,LMS���p(4"":��t���qjk֮���I\����}�X������m�А���Xߥ��	��%�����Eq�
��f�{������y�>�;�Z�}�P��-cU펮"���{������+�9�rrA@K8WkU��:�B y����(����;�<�r�/�����[8?T1�4xF����;ﳮ��/fpY�͛�T�a��_<*��4#a9��b�h��KNA�Lk4K���d����;L�mk���J�Ll�BR�J��!�����<� ������_�tU��Dۏ�[ȴ�� ����g��vmIuAny,=ÿ>�[X�$ ��X�"�q靿�A6OdG"v˨���؉'�o>=�ZfN0K�l"�w���_ߜ"�qc��Z#%���sMMM�؉8@��^c�A�}��a	����Wxo��X���y���F?O�嚘2�<u�� ������iL�C,�Pi,~��E%Mͬ�?�0fIec�w�60�����+�f4l%���}���;�x�>* �X42##��iixD֍!tx=mf~~�/r>5�"��wk�h���ы5&rkVAϗS�U��j��$k��J���H�i��*Q���Ǥ�ݽ�6	k�+-!..�@�gư��=?b\�Hh�0@�M1i0�C�m4�)$���u���fyw�j�Iֱ�uB��T���YYR��}?HD�@ �gHII-$  }O
��H=��{_��T m�'�ӓ���dG2y����;M��u3�ޙ��\�
����� ~5���4640rs�Dh��O��kN�f�e���Դ4oc�B����hz�Z���[\��*�~��	ķwU��_Vo�rp�m�,�O%���-��-FKV'�~
�ig���w��m_ ����
�����|�`h��s��Հv �{n��]����#��l8zm��r&�J���5����bb̝.�}oPw���!�=Y�bm�>�=��9=�OS"����^���;�s�A�����D�¡a`�Z����b��^�����k^Ȧf�O����aD2%}�I�Ym�yڪ��A��uE��ӌJ,�H�yj��S�A��ѱ��gΜ	�Q��g^�M!Zr�x� f^j�{�
pA�N��K�cv�^�y�ӎ=;�ݽ�GE�+l�۞2���������X��*#}d�u�f�#ݷӈ��Ys���%��]h�uP�֎��b����v{?�}�//Y��|��@�
�����[�op�|u�p�A�˾]�`��K�W�=��(�gw�ܴ�s\���E�T2t�G���|g�M�ruq=��TN�F]��a�u�� �������1c���(:n���(d���:y߽f~gy��ۄ�ⵁ�Z��݇��_�w7��AG`��y�jٺ���=�z��� D	zT�rW8�2���)$u��%}d��������%�@V�������}��=���R1��K����T;��
��0d������K"���m�J$A]���ɚ���y'ªЇ�rRA�^K��f�c�̖%���){�M�Y��Eմ�j�Q�}���2�""3_������m���v�Y�s�����ο����:F�Bf���˟X�yS��'�!���-j�/��|�UA�=;HxO�2�\;}M��$$W���A8�L�>�[Y��U�{~�̞���A@�K"�H��|�k�����14�3Rt�[!n3�[0��3���4>�'��6<�����W
}0S`D�0���l��A ϱm�}�D�A��PB����l���u
<���%m�9�����6��Z�����5�SL۔�V�Yd�HM�C-~��y�ٶX��ލ-�du:G�R*��T��H駉�e���u���TT�2d���?
��Ir�t	D��t���^d�O�מ\q^@�e����pj�#� pE�H#��(e��އ�Y�{h�2y�sD�׮�S�-�������?�����}CJ~;�D�&�y/$��^i
��Vr�cat���Nh�z���������y.��d�u		))��ҡ{�<Y,��p��悔YO� ���g��~�l(q�Xo�F�$%=gR�z�9��V�9!�����*0]����S�T�j5,�=I��l
�o3�\�{��x~���ڣ0�]��o#=�����<gu6�� q���n� ���P����V5O��W/T��?FkWX�Fh�5��Ci"�^����涶���7f����Pi����ga��[3>((��ۓ���fx�.<��wҋw��2��}����ӸD��r�������?�J����.�bhh�S�9`f���<uвV�G�!�����{a/��	�-��������|�kڕ�;�{Y`�+��Z�@������;�WJ�'>���ꗺ7��xoS�W���P��֣e&;��p����hh�o;Ґ��͹���`dY�D������g�\8 }	�i@�j���7t�f�=����G��?�ED�>�����^�+)6MYل���fz���0��2��h��B2mHLT7`�é�к]��J��_!O<A@w�E3�� :���t�T�h[!Ԭ~����>��_�&�w�Qc�y+��}��_�`�yWi�ܒ�Kga��{u��x,M���k���D��Z!]�|1�EJjCj����H��@����b�MŰ����1�K��V�Q���t����:q�q����Z�ɓ@�6��y>XX�����9q��{���A�6���i�KY�%�ƌ�Az���U�3(�w@�2;\Ѱ�gT����LI�������uO��F��� ubTN�3qe����}y6<��q��y:�� �99U(9����� �f�s"-����,+�����Q��*����G�f݊+xg<xQ��J�Ӎg��)BvN���C�����~苯��"����g��̼W����R8:� �����瞲`4t(��5	II�ػ�8 �cڢ���۞�f � %_ >AJBx,���`I�\F`'�}M�:��'|䩖M�7.9)i�'{�\�Y���n"�������r�϶����H��*�;K$��X�������|ܛB�i����$�S�9��0.^�v0I��s���O���dE!.}�b�f�e����L�����X�߿/��r�9:ޓ������N�*�Ff9���G�X'���-�r��Gs�@^��uuR7��Ǘ� ����>��t
��S���Z�8�]a �����⍂ܣ&��ȵ0)⤰h.�F1m�j�t�Nv��,�!P�}�������P�B^ю�牔T_�ǲ�������4t^=���ցu�PO���#�w���2&e ��Lz��J?/ Q��66��[M?~t��RӢ�n?IruS��r�7+��O��v�r��7!�aQ�P����r�� ch�z
��I�L�}�E�fu�	&-J����u�Z��9��ys1���Csmm��|ٟ{:v�)��˕��)O\y���]��ə���s��b%��Ӯ$/�h9��� %;��5|��<2%W�VD��G���x=op,���n�`��ޤ�w��{r��3gՠO�w�3�'���\]+�x&?�19:���^���o�\,���_�޶c��발u���1`z~����(�{���2�l�2)�bDD�[(
�����./!jVFv߿O�UⰢ]�3���%##+�[���o�6?y5+��yȷR���B�'��} �M6��g��X�m.��h�!���gN¿\���	OoV��.$!�(��T���
�T�����Mi+�-���[��JyD�g6YkWd=`���NS?I��/���.���n��q�y��o�<��g+p�!Rcy�૸c��C�?:�@IIiB*ɠ#-=NU�݊�g��?
�'E���`��̪9��t��^hxx�t,o�F�%``1F�ow OȨ�|���B�BQ�6Jn�N^>X�}Ǡ5^P�&Q�Ǵ^`��`��&��br{zEeeܛsT�{�7���
is��f��"�H�Gaj�����f��#��8�'^ v��Ы��8�j������+~���G�z��~������6�͗(Ҧdr�̨l�:��1��k!������0|�w�����y�\NA��U���6~&._����# ܺ�~�Π�_HV�}#����X`��AtZo9�r|��ʪ,'�{EEq�O�_�xO�m�r~�>pMX�g>���,w-[�Y���T��^�/�4�T� ���c	�˟��w �~����c��q�� d���Pآ"6��E�Qm([�������W�
ԣ��
�*37w�}o�Y�4t���vFww����b^��.b�'[����[⨦�O�>;
�L�ȍ=}�`���фY�f|�8z��ıxu���-C!�&$9 ��ex"��T�Q/%���K2,LI�󱈗I��+TAq�gC��F�a�Դ��Q���7�E3���}
(>>~Zd��c=��eW,wUm�� �ʿh_������i���o�5��}v��q�H]Ͳuk��X^D��¦�h�|wG�0Ԅ���ji�F��e*Ek�< ����B����9�zo;
�
���WH�u7��?�����/փ����%��^�s9b�y�%��bdsKU����"Sl3=�k%��݉�q�P@��o-������\��o8���^J�e'�@4�9�}����r}�m\aq�ݪ�Y�r$p(l�Y��\FQP��{z�kU��Z�� V��f����Q	k��i:3/)������֠%�9��Y<v��h`��3�$��2w�6P�Wyst]�tj�QIQ;U�kz7/���E�"�����:'���ڴcP����
M{�gu���7��&�O�z�rۦm�!Wl1h�g�}�nx�!>ǣi�F�2U{������Qvd�M<P�=}K�E���@[m��3���N
��r�-��,��<�"��v&���>�QJ�a�v�ٱ>ٿ��3S�"��|E��}f��F+��1J����ꖍh8�m�#��;d�x�`V��ϓ�o�={�����������U|�n)�%���=�����r;�|���=��܄Yvb����k4#��������B�����p�l�`8�1�3��R��dfeuk9�B]�n{�E�mph�[��C�#���U��k�P����� w���A���H�z���x�����i�+���82�X��{/<[�k�䊪���^��AL���[Bl�zX<c<���Js��l�%W>�I�,�����Y��TXcV�2Sq�c/�Ta�ꏗ��8�X���馄k@!>�.�4��aV���K9�ژ����4�J�3w�u&�X����A�	�m~8�q�uV#�>�W�Ng@@8=;�A9}#55*[��򇈥0��"����,����h%;s��<����l0~�+:Mkd=b~�P*o�.��(Ry�M�Z{Tl����?���A�wjy�{���Vb��F��g8�?"(È��qjĝ�����3�wF(�c�L'���/dW�M�����v�,����j
QRW7U 3�ߝKv��D?����b���ӓ!����F��2tf#�t��c�mUZ�rѢ��%_El]�^���A�D�(�����y�mԅ~��E�g/����*�Xk�n(��`���WaD	����٥�t0��g��iՠj�W��+��@��sEfs�Q`�121�6�A'�ܶ�әr*��@�y�;��9d�R�ØTv�V ��3�������tvPAee�Ƶks_��:������]7�uB��ļM{8��d�a�(M1��">�m���N�%�Y���f�e,�nN�ڹ�(�9�	����x��
��T��'�W���U��<�Յh:�j�-��x^<��.�s�tg*@��eU{FBF��Y��pf�$�3^@����^��� b��sw�g�Nݺӈ�������x*�t�+5myR�S̯�N��WZx���̽���y�C�̱�ǧ�2� �]�����1_NfY6DEZ�����/Ə������n��R�~�0�����J��e-�R��[G�z�噳E�~]���k+�n�qYw�N{�x廡]e7<z���r�0�V���s��rrr��u���'��(�&��~����������Eq���e���CGM�c�22`��+���,i����fo8�z��@�4��ొyyyj���P�2:	��0�uǧ�V��Y5366� �%�C��,Z�干�Z&p��:/�B���*h�8ԛ�`���?b���Hf�w���Iga�1\;3��D�����D]X��T��F$��m�it
�n��Q�r��򯹜���{�H�	���MfLdw�^	e�g��,f��uF�h�&�ߴ*e�.�d�;iY�qL^�,�	��ʇ?��;���.&��
���6���i�e�m!j��7���gBg��: �"��:Kw��E//�>�k�����d�-v��6�6jU�c����~d��i�*���P�|K��Na(��l"'�sE������xB�8R�˂ ;��r�?����8����Ž�݈�~?B]�������(��O�l����2�JgtZ�J9��Sv1��ĸ�?o��q�쩖��-TP���S�.�ﮁ��'��G���"18
�]����1e���E�ů�&L������S3����{��o�E_#K��!K��+Cͼt�; CDak?�Q���	���y�L�B�e�T��Yom�/���mPƉ -�N�3�������v�3[����(q��y�{��]##�����J���T2��?�#�>��F#�¦!�~�����#q��?~� +!�t��������B��QCC�Pp�ڿ�*:� �����hPW��#r:�V����R�Ą ���ze�cg�L �8r�E�?zp]���M$�p}��n^��1U���ì)��5_��	#�S^J��-���cqz1�ȋ+�Dp�Ա�W�g�S��'%=0��=5�#k��b��PA���緭���כU6$�H1�p�"�#��$����a,��>�-��]-�����qv���3,44#%��%�����*Vz yB��Y���I��ٔǥ�11��$���?B��ӛsX2Ν�%��_nH�?�")�^����K�;}��h2D�V��ͫlt�˰p�'��%��JK?[S��D%}z#����NZ 7�<ؒl�Eݱ�3az���\�ӝ�E|%/�nDF�����Zւ#.�<��o9�D������>�!$��)�-$���:�����A�m��p̆+� pl.1f�Q��Ѳj:�cj�^sbP��m-_��d���c���I�UO� ����� �O����;�Q�Q�7�a�����Oi�i	j��݅C5��b�e��^�B6�������/���K�ڇ�"�J�8�b|Z���!
؟GD�	�����l]*�-�򮤮�$�\E0X���~`��c�3�5E���Q��FF��[�A�go������;x��mvy��0��ʂ��;v��NB�rf�Rf1�O�^7a�ݻa��0Lㆢb��D#�UN�F���5L���d�2�"qS�T%ϷT�kj�q[f-nr?��FA��dD�\�W{޺�񚻟HZ$�j<�2�@�2�w�u�p,�õlXv�`8����{�'��A⨼cW|�3�P�m�"�����KiW|8�bm�4P�F>�P�-��5���^w0�܄��w�$�����Te��~��O�R��e+z8B�B+�m�\�)|�����Ȫl8�a�gs�fP�u�2�#�H/�҈����K�Υ�Q���zd�I��lO�E(�����A1��'|�|ES�?��Y�|f	������ʁ�@�fy5���[�m&[��s��M-��S�OY��
���� �Y�/!2_�X���_1r�+����hK�P?޳�9����]�u����.���E�O�^ 
�e���K�{��:���I��f��ajަ����o)�C(ڪ�Z�O��7���壋��+1��nCŹY�D�_�W�}l_U��+a��C�w�?'%=I��̦��FG��"8�4,&y	��]�%[�*���U7�-7*��Yv��`d�L���q����tHy;�"����"�.룳����y��*AN������=m��c{�$�>��]D+h��ƾkM�%��)M����']�/x�8P0H�p�1�#��V�ˎ��ԧ��}�>4�����f,W�+� ��=�_q���"��>�[�a��:=d�2�VR�q�-�z����F	��߶����Ҳy3j�j"w!I!j�n�L�9��√X��T�~�Ǘ�N�s��s=��G<���+��K[��d��s�Y�]��\�r��:.�	������8��:J��Ѿ֓�v@�HI���׌�8���Xs�X׳�:j_�{����ӌ9pSB*OϱB�����S0f����n(t����$;=�ɴ��������5�6.v.E��o �+jJ�������<o�b�Qh�.�uH���2j�A>B\F]���<QWW���_B��_��֐VҮ�!��a��f��fֹ#r$��w���G�hes��$%��8~�����?�1[��_g����<���K�$��ݳv�����&oS#8�+�(���i�9�w!k|����7츞\EN�9�[���M]J���V�J��Fu:��~��濛/��!�3�{ϑ薇����4����&u{�:�/���糸��X��3� �z�vS�"ch)��o�v���	�|�ʆ4���|����c]�I)�]f]>ї�\��J��KC��悚��.�<!!/*��������~��_d"t֊j Gj�3�N�l[�������D�	��f��߇�[����*���2��l�Wod��|gM�9W��<y���3����M�dm�-$D(�rϸ`s:����%j������[�؞'�\E��tՉŬ�͗1=%�U.�'��t�?�S����T�y�O�\a+)%}J���a���$��ܥFr�҆�v`�v�~�;�:md�}_a������������c�бI���4h����
��>/>��(���H�kW�TD�>��<���|AXUTx�v�����	���t��u �w28}����z��_�Վ+��cE�Ra��"��qG?�!o�^}�Y����/��Jv��Ӑ���x
��f��j�N$P�n8��zn��ϝa��}�W�;��!!c[ͨ��{��,	�{G7������pa/��>�a�ʷ�	�#�ȯ��;�엲��"�ll��Mca$�)!�kF9)�����>�fv�F;�khx0wM=,�����x?Yr������JEڹ�&V��]4����������4�c;���׎�R�y��%J���u��.-��]� 5�k���ڵ�;F����8����K=O����2 ��������<���!�c��^>L��Qํ��z��(}������*+�ه�/])r\�8��^|�RƯ��%>g�L��t�mt_�����˧�KW'r����ѕ�sZ���������d���wg`��͙0ܑ�Έ,�����O�4ٴ�Sm�N�b�u]�YnE3Lc���X	����ʪ�����:����"-2�8���t���zE�E��9��Zih��Rt��43�?�6 ����s��;Ǫ������H��Cޙ���{e��~]�k�'z�ϟ/�ڮ{��?-�V���;�;<ꚙ�@��Q�����u?��_��y�D21�Û�Y~Е�x���cu���:����uh���#���۴�p�r=����~�C���.a)��Y޵Nrs��ɞ�����c�����]��n�]��K��)Q��ق�\q]�� �i�3�%k���8���aWn!+�$BHk?@|��JK^��h�^���Jì�,Hc��/�+NAQ�&���Ƈ�o��_��4X���pZi�gk/��Ë����tp7�L��g�Q�N��G���%	�*/��3*��t�)F4rr,y�]�2
��$�=%6n�D0Ō�.֞V䖙��ۊ�q�=y79��5�����A�ϥr�v@�h	�ax�6�0cՀĉV���.hc��XF�f���q����OJ���:u�a���C�/CT�%�������#ʆxe_-�Xx�jmR�-t�$=�}��?��f*L8K�A P�ALFnj��yO�fl�� d���厾Y3u�2��@�E�,8s�VQ��_n"�V��N������HY��Q�W|�g#���_$�`Dv/7Ɵ�E�:9���&qY��ޚ�T֒�]���*$�ۇm8��rPo�(��<��B�VI�~�o,���:	�9.-u�Q���-���G{�IH����sj���ͳ��G��7A4��j8aKQ̯����s�x{��'$^���5C���QX�%��":�l���e�҃�ā ��Fߪ]�嵫�n�٥`-1X��N��GKk������>9V�6����2؋ʹ�%��pfc�:����8�����w��&����y�������)8��s���n������;61�߁{����fy��b�!�������v�#�0���q:�"���N�kԷLm�c���޸�K<z�+���0���w���~��?x��&���������u�2�f!%�n`�X����*��vgd��[��46�٪h�en��Q�ӽ��*�}~��?`��x������Ѩ�[Ȫ�PC	8�+QQ��fٱ��]J��+��ڎ_3J����%�#��}T�O�R9�7���gw#̕�y�2/�
���We�l�-�@�v�p9�Tg��>p'��ok��F|R��=)i����Ō5W��Mg͟>�Է��D��m��Ŭ����?�jG����T;���^LPm���r쐵��Y��:��{���
5��\��^`XWj�.��.L�����9UuN��^�i��^�p�oRRˌ��ր����$�P���Q���j�0}������6�K����NB�{`=N��7c�ɑZ�i�g�}�����st�Mt�o��BP96�?��+/�hi����VνKXQ�'�5"7l����LY
2%*��g%E�KXA;w#ĸ��QNʞQ���'�9�S���o�D�,���@��,T��f�k�1����J@0i�(b�����{�)�`Y���օ��^�B6Э�U֢�]0@�%&���u�[��5�z[ǂ/09�'X�-y4�N�5j���[�~��D,f�m�Be��L��J�Lt���Q�ۤ1�V�g��[����;�A��{�%�`��s�nɼ`r�BL@]J���A�T��Ҥb����̹� �	�O��%ݟ.Ss�i��3e��7�eZ}3MtKL�q��j��V���J-�9s���%SQ�L�=�`�YT�p{3����E+v�,D��:]�\�J}G쀏�,���W���wA0.��������
�Y��;~����x�˦cӥ��{+��6T���wkb��H��,��	�o^�+Ze��Y]f��;��O���1(%��Sj�_4�rP
�nB����a(�U�<����/�@e�B)�.?v�6Ĕ��ז����x�HImk�JW4���3��h�|��Ҋ��k��;�Ĺ�o�Vn$4&��ͦsw�E�w���+��^��az�p�/-zu����A�]@�oG� K����'jM����)CR��ܡ�{Z��n�"^�p���8�u�ͬ\�
,k�r~tm��SxloJ���R��馞im7L�x��Ș��K.��mK�?.:����!Rʙ�[&�ɇ�@��lի7���hŢc���q(L���S}ݥ�L�����:TN1tg�����.��U��D��%
r��s�QE
�D�O|��X�ɥ^�PGǼ�Se�ج���/G��X��}"�QՈ���6��iQ[�^�#�a:y%mfg�%���ف�\(�b�d�*-v-�k�Qz�}t]�=��#�"�AX��Ԁ�NӐk��U�:�rT��[����5�h�����qg/Qg��?�;A��/����j�����qhj(��ѩ��㼻5��@8�*��Y2�r��RHA^g`�QllF)�.�[��=�m/���-�,�B;��:*���a�d�6�z52��(�����7�-�ZLk�� �rH�8�-+�J^;Ǯ�r��L����~dZR��a[7�d�q�U���Y���n�l�5Ldb`j���L	I�!6,���5���[!)�
錬�˗�22v}�%���zZ�j��{_�e3�x��]��.5&(�##0�r��{)������)��,��g"��bn�!�-Q���5H���Qy�@�4x�e�R�B��*�D!�p�0��KU5��X9w��.�|>��A܃4�*Ǽ]"J��V�q���r��H�ti���9���f����L���3��~���G�}}}=��ݫ�7=W�͹�n>�N"`�^y[���*�fQ&�4���6iŽ��ȏ~txR>UN[�����Ft�O6��ē��Z6�Ǜw��W��f	0 ��.��3��Y��a��p�1A(������`*��>d����X�}|��׍k$䦈ې���S������ɑPA��T`g�T���p�|�u�T�U���=�Y'O�#ҀEqm|+��^# �贰� �y񨐤b��uT���:���:e���b+f�H-5�9�*zУ�P�:n��ˆ#+iD��f��K��.;0�.�S{�w�>#�;��'?*����ˎ�
��V�*t��F�0tm����k���&��4M&޽���qH'Ι��,]�1q�ػ�}T� �ͫ�j��	Q�x���Hm�R.5��k���d�FQ���|��<�>���h�w�jwO֘1W�s
�Ig<^� oٔo�2PtsO�&^�	�<}1h�8x�	��T4����#-�q��A����������Q�F`	����b��@������b��.�*+
���,�\���$��I͓�!X?�`�W*D��A'��Q�Z9��YO̿����`8���T��(��}ҋ����[F�K
NUڭ��&�O�~�;���MV~��턊����j���pYDA�ȡ��&@mzK�%%���HY{�s��`���lp�<F�~9�R$�{x�|�e�����'��]��9��ny���~��1Y�u�������RXz��j�o��^�P��&lyE]��>�D!����"���@&�C8�u����
���1Y�ʢ1�_����A���� ,2Ó'j,ꅲ���Ef/DD���{K�'�}�6��������q��@��WOA��M�E{�Jm���o��E*��rw~Ȇ!�+h8���U�n�Ssz��)�n�]Ē� @t�d��=p���,[�n΄��T�/�5�t�1@�/I&t�����Y�w4�}b9�/IG�PU`e��_��\���q�������Y��9ӡҵ��5���g�A8��ߧ�%8��Q�?;�I ��y}�;�ӻ���6���� 9g�M�� e��r� k�5��b��tP��ƅ�H0ϸ�;�_�dD�e,�Ӏu��*�����(v�FTIc�c�����,����0%K�\Cup�fkUc��/Kͳ�k�����iM���{`��CF���0������h/tLzl��E�%�>��oߞ�;�'}T��u_�s�Oꏡ;��t���,3�&۸�w/�t?3���b���{?k���V9�63\�^�:/����tI��$��,����ֽ?=���Rv	p93ĵU<�@_�/�� ��@P���:���ݻ�OW�� `s�}#�ݹ��.�}�i�� =�^��+'Ո�j����ּ�[X���q+��f {�o�,����B/���;~�L�k�7�U�p��o�>�~m؀�Ȫ1JE+�1ʀ|�����9������')�졽@M��;ޯ�{~�����`�T������h�������!�c���/Ϊ�n:O]0�]�|T�{R���s�"���P��[��Is��@�I�� ׀����o���q]�o�S��T�	[Y�ec�s]��v;�����d���0���-��T���x��u��F���{����nt�*-U�
l����������k����Z��_22*н�ר�X�m*�<���/�_A�t	�U��������U�߃�`Kb�*m�[����&����f�4_ٴ��IL����O�)ogWH����\,�J	<�e4x�z{����PU.���k]10E�A�� ��KA���@���.��H��r����o��w����]���13{?����~�N�og���\��˦�@�f_����Fjp){�$�iKG�@���%63RP[�E''���@_ߝ��5��� 9���n	����rF�}4t�0�����n0����P���5�*�R8���L����{r�H�I�:]�F�pX�8���K�y�{usYv�\�XE��7wy�f�\�K����S����V��l'����!<JF�����Y�Z�� �o.#�j�a��:���J�]''/(.f�������*j�7աF�P��xަ�֨CxH�Nf�l��Z�a��p�SQ~��ɒE�`o�4���T�|OFǙ���r+]({��͹w���/O��R�`^P�&�x*�۵s�P������c)åy��]�)JCK�S6Z�o�6�V2��q���IC�1��;j5�%��bUr��E���B)�/>�(M�#�w�R�Ҍ~|zQ��D�EFf@��\U�:U>����*�_u����F�+��2vpX|�R{jGк0\".=f��^;{��u>�K��JPq&��dčb#��m�|O[�Pp�Ҕ���^QI)"��I��Y�QX9�e��>Tv��,���LR��͊w��&�u�D���8.?�|�g9ǥ��Ҁu���h(��Î���m<kI�]R,��wޘWD�ݾ}�v�if�z���%�v�K�aG<�Ĝ�}��nS T,t��K�w�����d|j|[�P�ܴ?��ȫ+������ɵ.H��/�u�h�?i�jx���t\��-�������b��n�M���9�HԊn��������uaG?/:��v�(�0P����_���=�) ��_�Ǽ����=h���$s��'f�l� Q9�n,S�G��<Ixظf=V9��2��+ɧK�.�ՠ��44bɜgoAC��� ���?I�n�%��}4�1�$�Qc�n4�Y4������u���^}:��<]��)/"��#a3�=C��aO�s�۟��IA���4�D�.%�(���L�9�;gC���2���in��h ���I0k��ë._N�7����x��[m�	��m�6��7�)�k$�aU���,�Z���A�M��ű�9�'�^��l���֣�{��X�8y�矀��.G�H \!������&��%�o?�9��*ݩ���ڂHyddWW��*5�h��\�=I)�}����nA���t.X�ݭ:\��ׯ�MΞ=[�����$#���g�������+m���v�WP���y�N�J�(jc��1��WRP0���ඝ}kmcs�4Q��
��٤��A��[#6�W��[�i2D�(9�O՟&W��]?Ce,1�U�**T�I�ێ ���r�J���3�Z#M��k�y"V��ǡ.�?�N>}Q�s��,���a�	RS�t��Y��&ϖ�i������&�U�z����Ft��aU"�`���ʊ�s͔	a�V�o`��0�%3lcmͪ�t�msЀ����<�M_j�o�)�Gl:�~�A�$x�V���wp[�455�a�x �����	>�BQ{Y�Z��A{/��&��{ d���.1���E���]����Ll-��_�H+�Ԛ0�����f,---A�W���8~z$T���ux�_ �T�Ku![B�=��r�,**
���7�D���BktQO�:n��+�T}� ͽ3�_dԝ*
E��Y~��D��4K���%�a���%<,�U,,?s
��Ԣ���J��{*�nK3�O�:��P3(�>K�[[S�P�*@�BK^Eq�>$4�٫-�ѧ]UI�v��'�"��Ge�DDL���_@����s%���`ś���� ��[��fg�^~	B�te� ZQ_?j�Ay*g�_HP�RѬ��J��Ɖ����������t�9�-ͧwwD���-�z��`����7q6�c̻A�.�B	7�R?#�s�]��lM3HpS��������ϛ�pQ���7���M���cv�K4~��	2�������6�����JJ�G����.�ݤ�K��]x��gg�����mfK��Y��2����^����rB,ˌ��zA�6-�� �����_�<���\2��qE��L�MT� �C?��^��T�c�


���6�Y��K�x0叨��<���	��E]�al�$e��������"���Vz��W�+�(2S�*��,��Ϳ��̰����D����K��[��+�+Et33��Mᄄ���9��
�����?odZ0xeG%kk�͌'����]���pL{�a��I�E�8ېj-����qqy�9����ΤW�+�׃��ۢ�:�ۺ�rMq�޸�~q��SݢFq�F9W%	���R�gZq�#Q]�4	��RLŌ10� 4,E��ؕ�=rG$hV�n7��Y6`�$[���2���*3Q 1�A��1 ����M�~���u��������0N����!�LԚA�s��	�z m��2X���M=̠���Hu�:v���T�8N�Ee#}�J��l�[A%���j��$���!�VI�@^�>�-Y�8.H����WRJ���K��-��;~�B�QF�t9��=>\�Ѡ�JCBVXX��a�7�3;�WK��ʆ�b�+���;�E3뉽:;Zj��W�kvW�=4P�Rq�p���H^���,@ ��O�ulԺ�~#��mm�#ROjh�G�Y�W�q�Α�uL.��qv��A�����C���g�aI���{?I��]�AE+���B��	��񈕩��0�V�AEͱ{��� �gwf,�I���=�Xn ��>�C2�[�.We�xc�c-f����l�%�Ε/����� �|�r�W^�N�����c<,)�ڇ��1�f$nҹ��l�H�&qƚ����`�_:/���6(���l�s��B��el3����!!!X���;��^][c{��-���� he��y�.�V�5AA�k��-�O��.�H�����8>��R3���L��,MA���Ϣ;��l&���z{�s=9���M%aa�m�l�$����&A��fJ<�����i��^O 1&	�[��V��ȹ��"�fU�0���Y0�� v��Q��h���H�8H��N�~��$ ��u�� � T�<xd ǘ�9���^��\����'{fQ�B�k������TI���Q�#6�������V�s���XՔ��3,��G.m�Ti0��g߅��8�r�<���p\��;&�����z͙B�z�b��9��4���,Bk��Ȉ��C�HI��5�y�ﺽ�9����).���2m��qeu#���AW�xlg���)��&�i�v� ���@�Lsuu5��@�m��X�v����=�a>ݦ�;�tƷ�gB	��sJ��>�'��q�x�xk��o��a��hZ��IMM���g���Ƥ�F	"33s�6�(�y�:e��K�.�R�g�+�����>"�r@��9���˙��Zr�;���e���W��nҺ�&�6�6o�����rc���y�t[L����QJ��ظ�k�Ap=<�K�4���'�z)��q�,�K�k��_�:�%㸃�h�Wd1��%�Tv�|1��A��}��vV���S	�}g����x���ũфo�IN�t�?�j�w��9��� u�y�V0 E�gs
j�vk�@4U^
�����Z6�y6썐��b�\�onH��(w��xmS�X��IW�SU�- �`T���(�j� 8&�;�e���*�3��Fզ2$�,V�%E��β?Q��f;_����K>�MRG�L���y�5"�*���o�4>Y�QO:lf%1�j���+,��B)�\C����?�e�8ĕo���-��|��?�7��3��fb�QjfQ�44̿v3S�d�H=���>��#���P۵�9m~�`SM-ވuT7�>u�I��q$��]��2�f�H�����&R�9���(#��M� f�������Yę�<���R>J#��)r�'�_(�vE"�5�$IWD�m��*/�A�~Ri>粿Y������1
�V��A�/u=�5���9�xSч�g�[���[�	��63�v#(�
[T G�b���P]���ۮ��S+��W������;����Ԅ�����E���𰰰�o�+ܿ�J�������W-�1ϹOEW�*.�B�'��u�D�~z�+=x�����q0��{b�YYY�w�yY���_��X��HU��+)��JHӖSN�\�r�S�{-;���\I�~�y%�d!ܜʞ1�`@ zL։���^l%�kL:�c�Yσ5�}MnY5z�*���G__�;�ݻ�+L�]��8����Y��|l�/�S���.M�.Q�P�8��.<k387�
u�9q�	C�=X�cnd������ط���ːq��BQQ���eE���_���:̮��t�]��lu��(��?3���f�G���	>�SO����	�t>�R����Am[��K9W]�^��ư���[ۿ^x²,��}�cI��9)���,"��f˺����P�c���|yP��=�����t��	�w��e��*}��p+�}2����Y£_+*�|�SPxI��l��G���	|�jv���~��h����`Z�/K0�JI������J�����%</��r-��U��Yn�>�E" �������p����C�y�Me�lM.9B��c�1{�-{���vn��!I|�����݂��}�|э�M>�AC~�v 9��h��X��l�؍��^*rq�\�+��uHj=p�H���XMWTl�&�G!���g= �^}���@m+a���m�A�C���s)T�c��ǐ�;��rs��a��99�dk{�R9y��{� ��7f�Rd8�=�KPC �#�5/s��,���1��mM=����G��[�{<+iͬ�	����wzY�����Ge.#!�~�J�G:���2G
O�z��|=����|�u)�}fvvvSIo��y�L��� a��@�YH` Bvwwk�=�*H���tp�Q?����m���+a5��,���Yk�q	��V+��Ǆ.f��	>
�VR��>�P�8Y�CC���Y��Z#�Ѐ��G��Q���̑��Y�I2O�]W�N�i�@L�O�d�Z�"�{�n�������*�)�U��9���'?ζ[�x��c2����~QIL�
�/މ��j�s�H���D0j��Ć�NGp��LA���������rʴ��$�t�o���G�c�2��Dߵ-ܻ���_�����kw����{8��s�C�Z�b�d���ȗX�+�2�U����:��U@��xW�����$ָؕ�q��-��H�,�c57���˱L6���*����y�\kx&s|i �
6��Hkֻ3�G���g�K��ļ��wviӥ���o��N4l$��4�g��N��-��Xғ�*�?i����&,�N�u!}���y�A�c�Q���[��:a�;�2�s^7\�Fԛ���[;�n455!ɾ'�;�S�.$$�t��;3��p�	lV��/�f0�B������k�sۄ�5S���8�UAR�\@���t�7O�Lx
����L�A�,1C�v�!��o��> ���@��Y�d����2�c��x��C�~Կ�h�>(�糨�/mimE�=)!*S�(��3�7���`����n�����pw������.�n	ч���U�+�����8��b{?>&&'�7��_t8��a�$�3ye��ǔ~�'&&H`��Tփ@lwO��֨O>�����Bk;���ƈ�7�Z�{�gM��U`Z�a��r�gC��ˡ��E�3Q�P���j o�d�c��Q��HlA�ajN�C�S߸�:����[xܨ���;2����{����ƾ���J ����o�z��4y���j(w�@ɵ�O=a�:��O0k������x���S�T'���˿����K�#5�}A.��Z�/�:���<xػ���+�3�7/v
��C�����[#6�d�?�!��5��
�\��մ�'���
|{�£��LA���3���;�����L�CcAQ���.�伾R� +|�,�X�r���:퍋�I�nZ�C�d��D�)���ɟ�2���bpO�?�]�gſ��i� ',��Թ�� 2��o,���q�N�jK��8S� T+3���@+�v�WP%F=�@�)0��Gl^��/�ɤ�tWJ����n.-��<>.n�
�~t�؅"��	_J㦀k����g=vZ�	�	\���\L�4����A8�FV@@ ɀE�";�Pc��o����QW*�,�DR���L�vvյB5e�ƖLʣ488�� �P,�1�8u��l�AO�$�ƙ���9��Z�������������|]�?70��	��#��*n�(JųH����^=G���n
�+5�|F�)�|~;���|N�}li�h*JJ����)\����Y�ƽ��7�K<D#�����3�3�9��Q\��	���+�vKc�u���zl�-����_c~P'׊��G=�o�=��8�`��⣢���\��RJG�y��a�r�g5�D��<�p�cu��p���I��fC�N6����n�b�:VFL�+���O�5�b+�ѓ�@n}M>]�]��y�6��nB�hi��{��=����ۺ,�jaj;$lq���[��la��-�P�rT+�G�:��:KD�y��~{�b���2��_p���A�+2��=ٸ;�ع~�2>5�,F��Y&�v�F+����G'ܗ`w���Zթ��>�g���$z�6�>l�Y��������8 ��ww�)Qʻ;"��+#6pk9�]MV6	n�ö�(ײ�<8��/��rA�6^*Y��͋o�n���7��}{�d2��-"��1���-��C�F�	\~�;@�`gv�#��[P�ޠ#оjT<�M\1�c����/�'C��'hj��ammݛ&N�T��+iii����\�ߛP���Z4�9؍t�m���S�|��g-~�p�
nԀY�0�:����\��\�F�%g��"�A�0:�|'^2(_n�_�f�A�����z�ذ�[ �����S��ed�~3+�|�?����jO���H^�X�������������euyv�JJ�#��m���G{,�,���	)v��Cm<��O�Y3�����ϋ�M]===�v6�TZ��ja���RKMr0_�[���Ill�ZFn%�C���9�ëu����S����vj�����C���p	��5M����|���5OYsax�Qv{+H4X��T� �a����'��]���ź��Q!7���VC�Sj����Ѻ��1+�k�?��w��E���Q$�Oz�������wbk[��O����T�̰���d3+�l��e��1)�I������V[¨i��2P���5-�ꥦ]�͡&q_�b�|�E�m�kh.Q\��}(��K/�y#h{d}}�9|p���~��u�LlN�&¦ۙ�ɷ'��5c�W@~�u��j��n���窦�[��� X�^��q�	��&��#NۋE�}�_�t�-��Rz"�ϫ(Z�_�gXd�	f��+^�M	�.,�M���6�~lgg�ҁw�Ttߪo��0�Մ���+�=�"�g�I�ո��l��X�$g�|��\�DT�溹��qQ�����6mlCU
����'�>�f��j�����x����5�g�0�X�Z��@�H0Y`%����yZ5ƽ��I���phz
�A����%���eZ�(H�J�b`sv�=4w���S�ɜ���~��w�cs��a��o\��˂�v�@�wv��y�f�D���!l�徇"7�s#���[4��\���;���@��~����k	��7����}`�#��e�_5�u/3`�*6��p	 (�8EM�<��N�#|�Ԑ����tTT���Њ&����1�ȉ��r�2�97�Eoa^P �ϖ�j�\���e�	(��A��b6�����m)hi��2+	RMY*�y������<�W�"
�t8�:�9(sP0�n�7�y��R��iy�ہ(2wE�y�S����ᾯ��b�� ��Z7������Uk�뢰�����όﲗ��O�|`[X���m;{3�� `�!2�,�zM{A~~?��j@��W@f���8<��[nYB�(1TXX�۝��xP�Ɛ����P\#ȀTAQqD���䮉�C0`�L�e.[�.�%�x;7�k���p���063R�L7� �Cm��M���' ?n�K�a������J����\��Vg�!�>#�p��k�;`��hBZԦG㢅J��E���>��d�=��o�#ö���{�*~)�'E�����S�SO%��y}%&� j�����OMMq;.�(:x�������L HV���+A֬ B%��@F��pw����\�ŀAJ&E�s���#E�kk0��&�!+7W���q�֭
�0����w�< �b2�^(��~fa!3�Ƴ�:�M�����Ez�4�B	� KD���BL�7�6�<��X��L�yV/<����_��ݲ�<��Ld/�?���\��I����"da05�>�@�7�p؋��Z�q�@���~��:����}��Bݻ7.�$&
�<y2=��
�Oj*E�1qNy��I��_�n�@�3 ��:~��E�� 7����9)���%�^�笋�,8�<�KQ'Y�����M�E����C��� ��:1m>�(��p�lv�3��L��:*U�Yu6<̑�:�"@�N���Q�nM��������糹�S�cCZm�\�xr��iT�u#A�}�x�<x��G0q���v��e���x�E9�a���^!�;m��ߒ�W�y'��R?�EX� ;�A
x�?:R\]Xh���}%#m�i$c���[�'���ټV�-ޚ��c̡�c汓G��9#��!���N��	�����9�O��g�ARJ�X��#�$�H����]��]�i��I��v�ڵ2��Ω�	�i9�Ǳ��K�^x���.w)��]
�vJ鹯�	m	��j�pf�^ng�V����D����B��"������ᰝf�Usuj?̆��&���A8~�CE>oq�F{�z$��SA�Z�5�Z��3ka��uz^/�u�TK�S�uE2M'��g�E�� �y�s���:��9�.���
C�Bb�����?N�镱��E z��9��J��z-�����
BZ�� E���2B�MV��rIf�����?���3,6���9�CIlE��($���]���Gj6�"�$����2G*g�����Ka�?Lzd|)�����w�q"4����̩����-�.2=���2:6�4բ�}�I��(�t�N����8|��c�:��hl�Ŵ�#.D��%L1�[�ȋ���������~��s��U���ww=��qh>�#���ԏ%�⊤riw
�����/���MI�ew���z��c�^�|��g���{Jq�>�EU���该����%�$#;����fNZ�FJvN��Yj-*�B�H�����mOa���Ա=��O��#h�,��:*���#�!U���!�a�c��ڤ�`�ʌ(�1H��j{(韎<5o����������d�����J�ܦ�R��Ղ��%0�SW�[`�Y�Ӵ±��ܓ����������X���iի?��W�b.\�#����A/9�v���L�hu�꠳&���:��FS#�0aX� �9xr��������y=J�l�WN��w3z�p2o���K����ǰ���PwB�E����Bx�#Ms
�#�� &n��!Wk���}`��E��dJ��paݴ�
����+LZ�*y.��f�"r�]GƄ"d��r��YK᫼(��0��a��N�Յ�ss���[�ZHl�BP0�G���}K+z\A:>�0�G�8~x �T���e�%tx+��<��[�����^���	3':����E�*s'���8SAԄ#�y𲈦�w�D���!��G����ɕ���}��n�'� k�h�cEB㕡�Us6����G���$O� �R-|(�	�f�g�;!@�)㯼$�rPp���)�]���̤���g�|4ӫ����}���*���?��yɩ$�7�x�w���(r�����p�`G�o�d�������Iwd<)���ǘl�&=��yìTc�}*�uN�
��e$.�0`��9}��눧2���S꫹sW�0c�`��������������49��i� n~t�4U��	���[�|���?�A�q���Q�dz�M x�&���e�V5)q��pljݝ𳢡��'=��o��8��}�gḣL~�m���9C�ݥMBH2:�y�{=�	��K8���y麉�D�=�4TIP��=�m��o���N��E\��
+5O��j���M?� �2X�3�G=�S�^�Z�?���xtRfǦ���G��S���Hhx��;�����|� 8����E�b~}s{-�M��i��9aǵc��}-[>S!�?_|>�����0A1��홁IQTM�u�QXm;2����.ܼ�RO�W�!���	�I��R���7�'G�A���1��Н.krjV�����OK�*:?����	�`K1��Ç4�^�k����>}<�����7,z0g2��5;[�+=;+����ɝ \�Lv�g���c�gv�ޱ�|?���ĐF,�׭��P�.���c%�b������9�-�F$̀x�-�P��G���T�+?�P���Q��B$[����i#�dEN����q� �o�j|k����VD]��:�jh�n����������P�$x�F<%j�A�_�L���@�A������`\C��hp���E>O�LIX)�uppձf5=],�t8��ZC1<���^Q��c����V��:BJ�d��p{�)�K�-�l$E\$!6��5wUҏ�i���n�"6_3|<�hr����Hk�{i�S��=B���L!ըq��5Q9Y�a��Jmk	"������"���b�ݦrJ���>e߂�/j+��gK^� g�@�9&;�Z~.��PH���=)).ﯔ����U�=��9� \����=�hOǕ�����'*��q�M�Hlw��G�2`rD��q�8����	J�Ft���v>������������2��޾~��|�k���8lW�X}̌<��fw���
����!��$>j>��Wӝ*?�����9�Ga7�/��缁6��!��(~|6bXq܇^����!��(U�J�n��<h:���#~��'�̚�$k��I��OF���"�բZV�^:���h��]���y��n��P��~��ˬ7�=�/��G^�^���N����cʭ0�����m�i�0�WJ�s�����x�P3� ]Z�ۀ�;����s,�$��?0 ����rʻ��<�W�w�[��=L������P�U� �,���"�sW|�P�[�s6�V�@�>
z2��(e���� �J#߹���~���3��?Lk��o�l���׎��W�{�+��&-;�)��t��?b����ō�đem�w.D*g%~ǽ
.kYζ�	����Ը^o(쟍A>��i����`���������H��0�Xѻ�&/[���ԧT7ʰ��Ci!���/c�v�gV[%a����#��-�࣪ߚ�p�P%���+#�dE�m������ҍ��W�w?�`O��-�&P�z
�|A�n\ߖACߨ83�=6|ê�M&#���g`�����l��Q��!�r�V�a&E����VB�c�hm���rΟ��vs1�-s�����~Xd�K��Ƙ��2F�݀�����u�.>6�����#L���6֏�6O�\�u8{�փB+�7�]����?���Z�F�A�QݘF�4a�ۤ׾�x
Tz�=L:��������j�����33�/��z,^C>�'w7�/-��,����(���'���ms�T�n�:�v#T5'�xb���ǚx2�aw��GQҘH=n��+�;�
f��N�Z��Vm>�ȱ<ˏR9_�,�ώ���m��W��"�(�S���]���f��Q��/8�F[�N�J�vR�����wq�]U�����^9���s������K�sI3���x����h?��E%�4�JP֚�G﶐,r�z`��'��5%��Π#z�D���-\�����p��X�F0�%�;�&ňز�FMSo�}�~�� A8���$ӟ��V�e�"+$���7o���6W�����_�o����J��R��U#_���£��m��{y��f��*�XXF�x[5�8w�	%)��Z��'.dN�Gg�E��eu���|n�{��%���ǎk����{�Q�lB�j㷮Y�vͲ��e�׽|��ó�X����/�-��w���Fje�T����H���J����S+�[�;�E����wS/�O�5��5$�z��F{k�͒��*A3��)Յ���3J��,ײ�c̸�4 F�'��o�V���s8oV+؁���FlÖ��5�4�u	ڵ�O�qF�c����ro��^!T>���tR���P�G͘�OY���d��"�����R}�s	;Uc�l��Sdf�"�`���ʙ��U��"0D^���2i��ҶN�ѐî�5��e�:?8����-�[�X_��tW0c_��]����jQ�z�o�+�M��]9��±�U2���3U�_փ.{<O۰Ê�&��^v�]d��.)RB���[�i�z����
(c����R\�1�]c��f}{罘��4��9:;�Ze����\�i�ωA�M�u/mZm����r{��g��
���Y ���CF˙���H��M�ޕ���'��k?�'��IKԫ7��=L�`�+��KV��F$�u?�^"�[�e�>���W��{�yw9�Q�˘3)��эig��~t@{3+::tʎҁ�j��=u?�iw�ʾ����ݼ_��טH9q�K۫%���|�� �3������w����+�2?R���=�K��&����ح+^j�X����._9=�b-8X�������_��t��J��ثsQ�@�j�[���$ݭJ.D��=4�!�^W��u����?gf�;�zl�u��h�$�Wd��M*��z�?� �o�Þ�|E;>�}y�l��G�R��e'�u�M }��	4k��G7$:���"�h�"4��8�4{1�9�J���>������������=����V�_�:��v�"����rik�X;f���Ĵ�P$)GHu���5��2�%�|Ɍ;a��|N&#v]x�ŸLci	�-��jc��4��(��mQkt�eOd��u��`��J��7�_4�;l_g�;�b����Ou�?���V7"y�v�����.�t��ϊ�&�8����y$;$y��Y��h�:������D*-����s�-�8��W�=V��_����x�0�C�Ϣ�u��Qn��I��<S/�2P�A�����&�|X�K��hb�y�V���!������l�+�*Y�����%X9{y������5�X�Z�-�kuZ뤼�m�V�룻�_^�q#��>�.vf_�<)��ƚK.d��'�/e����knu�Y'�9PT��31ȓSU�{��\ C=^�b�z����İOl�ہ��2�<J�]�_�Om�����h�O" ��u)���9�UO%�g��^��f�֧�ܼ�_#	`A��E�I7e���Ͷn�oفirU"Ɠ`������H0�V��i�Q��'�,��c~�����=�S-ϸ/�u_ko��d7v+�(s{��
�w5×\��Rϥ��a+d��{�����}�YU��/3��Ņ���3d	���-qɮ����*��3N���s	9��ӄ�vY���uA�K`I��B|`���7�{�����|��hR(�f��qQ�"���}b?p1Ew��X��n��VZ������̛���#x ��]l�FN�	-�xn�w���Hݸ�ߪ���PA5"m�=�2<�և_�^Y�u~&��K�9�O�����=�F�@ �g�Q}~���l�5�����]G�O�͠�>�&��;�x�A..�֯���V��o�hH�e Η�k٬��?��9Q0�Z��?W�r�E�;}U�[�ܵ��F��r_�G֌���7ս����!m�X��C��� M
��ۯڝ6@c�\�k�؏���v���ە�>6����RN���7��5H&;���+#y-r`Qi8;~��P=�����qP]��}n(�M���o���L>�.��R�}���<�[R��T��m��ҖL�dP���mp�K��]�.�vU��WLb��b6#秹�߱.*6D��lƍP�0�ʕ��i��� ne���r�l�����J���y����nm��7jl�/��O����U�=�$lV�N�}�j����m�����[����&�[	ඞ�~Gw��DM����l��~L;�V���6�s1S��v	d_d43��Oo:<d��7����-�*�{QH���w�~���O�$����C��k��FD�r�݂��+��LY���,$>ckܷ�ګDe�1͑7J�R�rDdʪ*��㯓����5׮��|Д{Ҩ��W-�NjJ�&щ��WFF������,6��ug�x��1���F.P����m���Zn��Z����es'd	�$È�w@��PF�����m����9��*�����d�����W:r^���iۥ��+z[JӮk�h��Ӑ�ok��< ��1�@����$o��zF°y0�0ũ��C��p`�R"�4�'hN>���g>������z���ԋy�M=
`���#�����.�y�������$KIS�4TSOn�k_(1}��J��U,/�t���]joX�EcquK\E���]���%���	���.�#l�s�(�ͳ��W��hBh�SJCS�-t��i��B�g���nѽX�j~����WC?���5c3�e���bоv�B�#���$?W��Tto�{�uE�K�,��r
�~�P��Q�?��DT`�m�UVz C
�کW�`j�q�QJ��Cs7�I~%n��*!����.e�Nx���p42\���k����)��"���iF�{j~��=�2�;�.s����Fd��5�;-'��t[r��-ɯ]�w����'��"k�DY	��z'�n�n��S/�71��`�X�CV[Ս���,Ҽ️!i���N˧��V��|��lK�3���\tC$�Uv�q&ԛ���2G��?Ao���[�ߗ�{�Pl��O���E�^dv��G{��XX�R$}��LOn7��Fg#�h+!'c̷.3���_���d7����T�c�D���+�kP;��ҟV����^k2o]�^���)-ns} �?��/��8"q���Fó�M��ڼ�N�G�e���ȧ�-phJ~/���1���^v�f���mL�<%�@z�_�9���P�`3�)��Y�A��B`�n}Ê�6/YY��Z�L�D�M�c�G���5�J	�0;�]�1jw,̥�d��F\m����a���?�!	�6�k]�m7�7-?![����b�i��DK>��?1σ�����G�e���o(���&�<f��W�ϟ7��ߍjf2+�d�s�4�I7J+�moxhUP�o��	��#�}m.Ĕ�>f%�����Uu�%�T�h�_{$?L������=�.������b�n�Y�e���N'��,���٬Rǟ��0�9��_7^�*�)7�[p�eaAΟ%���K�rɐ��)�b�3 �}���#g���[�֥P����$�RPM��r�c&x��KU�ʥ���~��.�n֘C����`Ԍ$���q4w�G&{SO��7`XD��>X�68��e�S�<BWC3�Q�B놋�)��� �kD���iܶ���
�V�q<���+� ��������R��#U�1�%�c�9��-d��QywO&L�9e�xJf�G.��{g����+�Z�U��ׁG�̮�~�or�����9�ػ��0����=�f?�mH�<��R5�����w�6Hq>�F_�b�_HǼpD�9 ;�X)y�#iQ��2���F��X)#��=��	�.��;UT�Ei	����<�]�S7�ւ�*��2M��W�&�`n�TK{��8[��E/�~#2�9F���J(n�0?�u��5-����'�|o9������酧���s'��k�3�,���>0�g��3�.�o+��<��H���}��M���6>��1��/� ����C��j�O�Ed�l�����UK�uQ�n�������oR�gf�3��H��/HJ�y������;,��3Ԣ��;p	)[A=�CkBn�}��O\���\7��ƖS������m웶*�� �6����������܄�X��n1�Y�.u�߸ԥ)r��6��O�W�~�� *��k"��h"8(Z�wPr��JP+&(��(�d��'Xm�� Q�0�n/��D�����jcD���2WcM�r�z|@��w��io,xu�N��ҳ��NY�v� ?���g ���"�Z"Θ��]NZ5�����uܠY{�ў��[����;�O��St�4�s}��ܪ�G��:��:42�{��.�ݍX�?��g���^�\奈ˀ������3Y������zY���J=Ƿ||�떽�s<v"�
�� <�֤#~O��JT�/�����"6nV��UF�B��\�?j��[�Y\��UX�iЗ�	N�~�/������f��{�ڴ�5�����Ǵ��mOm�/({��8��%��x{��P�}��$��w���\�22�Z��X7��=GIM�G����hv���b?%�j�_}}G�i��j���ݥ�������kBq�r�:��oBF��R>IFشv�*rǛ�]BY,M����ؕ-�$F}�����`���(�\<�ܘG��G{qiY��{��Ve��|��۝g��n,��ys��8u�����F�S���͠���ihl^�(�t�H�MJn�t�ƶ~�/*0勫yuhd�b�ۥM��;4/����bg�_�V����nH�� ���7�¬�|�,'Ä�	/�RS6#�NS{��ot�ě^,i�?�g�&"�i�#����"u ������-�oc�dԻ{�3��������gN/\*s[.�NI�&�g�tgEDyL~]�x���� ���|��U�e,\�Y�p�eR���o���]7M"�:;Q	��ޝ�Ӡ�:{Ũ��� �횏�k�7ʴcm3��t��p�1��s���6\�| s�Cw���:.W�3�)f׊�N�y��f�p`��t�"�ؿ<�yku�L8�a/V
�(���o+��EVy�������\S%Z�+��B��h(�����|�&R�J����S����J[��Vtyk�c�#/C����R��򋊳�������f���H8|����09��i���~z\����刻Pi��V8����vT�����>�ZJ_<jf|2[����G���;�'�"-��Wq��Pq"ߜ���e2�K�>~��A��*�H��,��,�����[\/�y�Ѻ�����������R����8m�Yy�������#Ӵ���b*8��-|s}��A�~�?v�ց��-��Q����o�����L:kU��_v�\i<�<�b�:����1!�����~F�f�Zi��8ƕ�`�j+p��ۙ8�5���%�xd���}�z{{͏��F&�q'2rU8�ߏ�?�7xU�R��([�//��X�fV^Ah:䎪������9��w���c��^äѤ� ���~pPu�;��[���{=��/������!E�Ǖ�����E����,Rw95���DsU�B��B�3?n�H=��bd<*�UCI�����:+�=�4���2\Yu-�3q�m;a��	.�[I�������<�f�����2��3Sk�w���G�3�/ ��à}I�M�����x����)������K%��FdƭPII��$[L����Uv��e_B���(kSc_3��:�c��9}�m|=�z�9��~-����~�^'/jj�x0O��`�Y&��E�"'�m<�͊WK{[����ZY���Zr�eד�Ξ�f�)E#��s��Ӂ"�?|�w qp8�P�<m��<�/0�G����k����]ΊFؽZmPR�^�������	�+[�|��A�Vk2�ɜ���S�+ݢ��j;׭�d�Ю��'P��@�w|t�l�� �v� +b��_���	+���Ye��S_Y�eWz
*��$����_@r�1m܇p���/6rP�{��]Z�d0��:��J:eQ��s6��m�x8q�?��gf�b���g�ˡ�x�ϥ��O�B>(q��H3�DAIk��K����߽M�J��ge�7��Y�W;��f�@���>��*��k0�hefsvݏ@��CU>�6�>�5�g=��c�;T5����F�a��~N�ܫ�*�6��yx9g5�Wy�9n�6�R��\P��պi�ܿ�.D��J��m��hA2{Q@�Or29��`�Od��~�DE�ȗ��xxh(��DR0;o�E?�c�:]�V6�ｌT`a�����5��N���9j��_�nUߵ�9��yvBO%���ߗ����?�M��QDR�\���# ?�F�(�餒nj�C��c|3��ź]@�����H�o]o�V7��$W��P6ϵ��� a�f2��OG���ǹv��ח����'NK�˛�x�o����^�C4����[����>�gm���S����B�o��I���2�Q�ވw��3U�ϗ���
+��J�<ڭo1i���,��$"w-T�HU�������	���Xg�U�B �6������<��\�b �Y�=n�!���P9��Dg�V����.�5ȱ�����A���|c��~ab}^WH���yo�i�T�$-��gy#m����v�1^N���Ku���(q��y�좘���P���l���Dd}jj�[�ֺ�� ���J�x�b�d˫ ÏS�w���G
Գ,s��Nw�����dIξ����f�<:s��zk���t�J��d�;C`�t޷}���XU'	��m��Ʒ��T�O<	!���y��<kF�l���o�n�$� 'O�X��N�{��Ȑ�v��,����U��D_���&nњ�CZ��p۴��/�dP�`�����=}�q;�+�p䫠v��2zgm��+��0`Oi�ܓ��`�O|�GӒIZ<AE�&P[Y��;�]��/]��	L��4����okȘ~�
�!�d��ݿ�"-}h�6�D���"��I���%e/��5����/\_n=!@K��m^\�X+�s�6Y�GZZZ�Բ��3������{_������Z"�"gfvޟ����4P���w<21�J��v��=f�r��K��o,�Ϝ�{O��t3]x�������v��{ۯ��<�'i=Ruy�>s7xm��Y�R#ױ���4�J�y��$p�J�3;oD~��]�"5�Ɩ��A�([�bf�'S��N3Ή�cc�F�r�o��]Ui;A��Yk�Ϯ6D־�C���<$gо�����;��̕+�B޹�d.H"�d��n�w����,�f�o���O����c���@Q&�*"
{YFkQ�bo�s�b���'�W�3#�����oh�]��P���H�ߔ�<��{��B�"�Y�����r�nTW�y~�qr�4�#[�pg��mt1k�1iϕD���'���O ���HW��uWܧw����b:��<�9��JIߜ�k� ���H~fH|���}S%�Stg/�m�>Q�	�h^D�s�~�.���@�u��ՄOϷ�4}�5�R�~M\��dp>؛%Bt�T��<7�j��V	r,��J���
�uo�!Iμ
t��@��h�.\�3����!�����L��B\��$�f�4I�[x}��B�{�\� _���WEUV����g�-��:��jJd�qc�!��c�X+3���������)|�G����/[�ͷ��qp�nA����\+��NG)�����i竀����v�'��
��=K/TOܼY3e����'k����%��)�nR�G�+{U�ʯ��PyY�R^��(2�rX�Eۿ���'at�'�]X]�
���X�
:�\d�;���{)��1�D B�9Q;Y�߸2j׶���G�*��3p���&�3sm��睛WdMo�`�me�-'D�� *�\�;���������5r��1?��#�ٴ�v�����܌-��a1q���M��}O��m�����bWd��S�u{�G����B(��� zN�2��dĥ.�"���f:v����.�ο`������j��T��	(���Uầx�G^��<z��ޝғ�tKx�&/ѫ)E�����m�U;@Mf���m:�E�o0�������B �͕uw��b7�`*�F���W���6�N5?��P��#5�uKV��i�"`q��d���� Vq*`������JI �Qvk�$�>ڒ�%VN-���R�^�_��Y-�O���]ߢP���������+k��F1�`vkֽo/KK/W�Y����Z��[8]k��6{M�VbF|l��zJ���l� ������!Y� �fr�S�x,f�U:&T�Sעuv7�b���(gƩ���TOk��]�)�ڹvt���N�1���	�\8w��Kƍ����ȓ Oċ�=ri4rp��Q0t؏Ji'��ИǮ_��
6��'k ��*���u\&���0�Q�s��
gW�[�г�B�"өyHs�5�9:�3,��qXOMQt�faT~�6�j��[�:���W�E^yݣ�@no�`����J>^��>�pO����'8-W��=k��>��;~���D"��|���%Y���&�����Er���^b�}�T�d�e�~��V��J[zwu-�e���8���qxl�_9^@��-A@LK@��l*DUKZg��MI�|�`���$��x���Ċ1�H����|%���4WA�5���p0����"�⼳Ra�n��w�u�;��:�r���L�*�a�?V������k���~
�P~�G�gU��LG5�_m��b%>�\CS��`P4��gP��i/	������_,�Qt��){�i�1pM��>�9���v�ĉQ]�E�<���-="}��dM���w$F�Z�,3�s���J��8��'�zm�`�VxQ��ʫ	
,?���>�ih0b`���Q�9�!�p��!�'�u���Xu�;
��ά�ҋ��l���� 1B��~jgV�!ndn'�,p_�t��HC
w �җ��TF|.bjW��ʣ�_/.������-y�=Նp�c�� ��[<��̾����Оw�,u$���e 1��չL~[���b��o��"lVg�ܓB^��'�_�H{�{�+���`n��}ҍ�8���-}��-�&}��x�F=�\�7���gf�E�K�϶�5�@W*�^��睂Ʋ�����f�S;�l���< ���5� �{ t�-?tH�]כō�$h7�ե�R-pߜ�S'��_���o.o�=ڲNQ���S�����b���A,{U�`�$kOt�y�_F�l&�rs�kD�d���Q�(#\�� :�)���A:�(W��D:oY���ib��.b���M�����D;5�]��7"�����g�sȍ�\Cn���ݶ������+��.�S_�Q��m��s�R�vA�a�s��wJJ�}����e\��琝A������-�7ߐ. ���btv��Nu�)>�A�%��}�O���^�!�Z��D��`������?zԎ-L\�l�cv�Q~�qr��ę��^��H�()�� �|ud?`��7��Vy@9����r�H�8?��eVmY����RD��"���!�Y��*���A�d t�|�b������<�������Ǽ�"��d:���`~q�-����?u�fÒH��r��\��2�Ā{�4���p���Z�M���FT�����H��m�0ˬU�BڻE��C�y�+8�J�(ѳ��~�U=����C��ץUUvn�^O��s�'yU�c�����{n�w����� V���y�u���1�3���1	3R�܉r���f.�q��c�_/�W~���<�z�S�r���,p�%�����끿"Īx>�o�)z���~�(�r�86jo`���6�4@Zth`k%n��(H�d��,��B�)��M�9L��,@��F�Q��)�`����t��gZp` G�D9��kr���q���H��%�Ȇ)hƻ�$�){}��`�q�y��[�r���<N\j��3�#7���ж�!��W��x=I��s�DxJ�D8H|h~�,`���pIg?��ʛW({	����ʠ�)j��m�&B%w�<��D5�'q0}m��r?�Ζ]�I��\�O�I�K5��4D��2��:��ʍPHne;���c����d�ߙl�/�;"[y�]��^��L��f+��}q���_�/`��$y���=o&��xmh�/d�X�������G�N�9K�	�|;]C`9���Yb\��,�*Gʠw��9�B,�^��+������o�W�C��8@�=���(&Ӏ��4�[�祻̄M�'TC�h.u+�v1It��2���Qm渵�~������
�l@�N�䨍�����������l��.��嶝-$�(ՠ�E�뒡6R��>��g"a"gxL�:�"B��.�)�Y����/ݠ���ZO��E�:D��UH	��?�K_���C>�=b�W�CC��`�(1��>N�.F)y���	�aǱ���͙΄�\1�d\1<��?����,�gj^Wùf2<{v�n��s`�c�"�x%�`>� J�������!�s����;�T�&z'������?yu7�s���e ;���^P�
�	��k���>��x�V�j���# I����Ho��Q�/Sh��|sA�9F��PS����&)��O�J|����/��b�K�ڂgc}%7Ϯ�֎B;��j6JfY�o�m������4���0�d���r���.n����ܚ�RŮ�e���L���n���L�n����X�]��F^zi�>Mr�<�k���'��7�>au�Ǿ7��p' �D-��C�׼���qG��?⋞�����Z[�//k^�/5\O�7�����J��Ǉ=-�<&;*���g�]��F�H���;�n����'g(�!�G�e1��Q��/҆8H�M�.���շ��ZY���O�����iv�<�oK�� �}WZ��E��q�	@�����1��@OLH� �·�.�u����)�hB��E��Ѐ��x�#^��~J�4���n��ه���� ߮-���s���$��a�i=W,ds�����u��������t}��$z�(	�3�`�Z��g^�����7G�RJ>_��؛�|�58ٗ�%�$sY���A����"�	��-��[6lKy|XLL�<G�S�c�Z�O=&�Kx<�(���L+K�}b�j�h>D��|<��Re��Np!AmFlR|����z�.gW�,ul�2ɪ7[�B 9�X/���p�D�'��]�G)d;Hٸ������&l�� b��瀚+�����uU�]�T�ߪ��_�E���E���$U_�W�0�s�t���x�����+gj�n�o�˧G�������,�i��J��ܸ�%������i�h�~X�&�A|�����[��}��N���W~�̎$�.\ƙ�X%4[�p�/�e��7���}�O� ��]�d���C��2��%#-]��u���I3�����s��eŖEm/��(��t�i��q�N���0BUO����f2�+<Mz��IvI���< k��A쵈[_�|d�pugc�pu�o�0������z�ŻP�1Y�M�k��nص�L�z.G�ua�� �z	����:'�����J�n^V��g���S�.E*t�MX�'����f�;`z��;m�-�EFmH���g��)��Ë�q��ݥ�+�Y*Ȫ�/�@�˿i��
E�V�6ͻV�O��!#N�*�']��[$�l�2��t�ĳ�v`GY8�f�-m6 N�4���Ch��;�3�z�8>�p1P������t�-FC�h��H����fv'tF|���f$��[�0q�jY�u6%�k��G�!Y7v䶢:���T���i�\��H]�!����}
�m-��l^���xm
�����*�rK�¨ۇG�H������ڜy�5��ܘZ����&�X�lb��9�/9�/�T����~�^���Y�}gIm��̡κ�B�y���㟫���9B�bX�a���1=!g(oJ\ .Dy\0)�����_��u#�a ��ο�W�
Ű�y���9w�`mR�[vd�i7�������0�CK祦m}|O�Tl�p6rr�(�8�E�
I8�����1��~�TyYk64�/���=r}�躁+v�W�<��Ũ���N�g�m�3�Yz�Q�E���FO��6�	+�MH���Rh���g�pB�"Q�E���j��/�u��3����v=K�,95?��ɜ��Zㅨp�#O�d��bF0�/����i���%t�֛������_�x��[�'��_�ލ��Ŧ��&��"�?ȥx��N=���f����B�$��wׇ\���(�_��p�WD���OB���t�ǱO!��-�pN�ھp�L�a�pb�ۅK��W�ˬ��,G����\w�$��{���D2c�ĩ	�ΰ���@�W��_\ۛ�{���q� ��Y�a�I`T;��c�����U�)#�=5Bsz��,�����,M0U38F�3�Iv����4�_<n��ϔ��<mnk�g�����	�M|_�YG���U#hn��R�6׳	��^ÚN��WJ�����Z��s����N�QY�~vd�z�{���&3`=�o�6�4��	l��'��� ո�ee}@=yQrAT"ڭ��2�Yk�4ۧ���a�VO;#��F�\8�_A'C9�]�~��������0����Gz2uZ��.[�.��Ns���f�Ȋ�w�������Y/"���������숺���L�{ Gɏy2	�`�G'7S(�֕�q�|&X./y��M�s 7�+�_����&�Ѕ��U��-�M�h��9	j��x��bt�v8�b��ฌ��ɷT��5���W��ή�������q�x��#z8�͕�M��j|�woL��lEK7�i��͌���],�}�˕��[7�zݣP�ܘ�����o�������`��5%2�`Q�b��۹y(���Z8r���0�?ZG��\�j5����(���ICW�%@uV����7ä$���%���`� mX��mE]-��p�$�'���Ǳ�U��XO�O�v�N�z|�B9�QM�	߽�}���C1��}zY������ھ�ע��ֆ���#~�\O���&�ͧ�v��������:�T�7�>;3*�������G��e��Ps:Pf�aP�U�F���Pv����j��D�V�4���7[���t��35�"�.���W^TIU�+C�<(�5����F	����qw�1�ƲK��S�e��Ү	\��������_��M�O�G4J�����U�m�L� bi�v5�I'o���·��4�c xZ|�6�%]��o��ՃnND�g�zɖ�a��k�uh�������z��m����i����]D`��ۮ��X���F�`�r�NA�h9a����>$�jcq��ʺ|��GX9���c��t�#�� �>a�g��72^��/�JJ=ڃX`|]��6�:-!���W��r!��e쟹�`�����t���\S3�ВZ{�D�Ͳ�ő����_m�\B�~�p���N�7�:��U������cR���R���9�zf�̫fS�t�."�wZ�)��.�5oeG�7�E�=�E��^��=�X�C��q{#g�j�X}��@���R|�5T*ST����������?�;�0�E�����e��h�����7=��yq�����¾�wm]9�`֣�㯥��5�?�[�".���0��8(��RU������W���h_	@�,IUa����^k×�6#����~�N�{�.���)�g��_�7��V��a�7��|-m�v]��Mh�BK}w���.�������of�c �Z�aS{q=6^���$���h�@/�]����k�6>���pE�BQv��9��#��]Hӡ���jr}j�5BK���J{y���c���Q-��ɰY���:i0��%��hN���xaU�+����� �v�����H�� }c������H�ڵ�:b�h�֛���R�z��L6��Np�f��ADu3�������v�g�)��R��������;�(9��vO$2[����55�x�腞�h�,�:Ũ�d��_q%_F�Z/� ����i�xmd��2�Z��n�r6��fQ�����,v�kk>��_�ߝ9~��?���l�ו(@�K��W��w�s_H��3}��3g�ǩ�=x<Wڋ]�<�煟���O���#�5c&�H�Ywc��a�	n)Ξ�ݔ�=}Xw���ag� �j"��6���J�#�-m���:q'�ͯA{��u�M"�`c�;�Z�����M��;��Ѣ���~$o��<��2��ݑ,y�n���`sf:�eE�j�9�����7�nN؅\��ж���,W*+��6U.�ˬZ-;y����B�W�,Zh#��_��o�4pȈ�l�Iv\�U��k�7�1k�/%]���EW��T%!��F����d���]!S��{�f&$�Z]�쳡���~�D�_�leIp�%��Q��X-;Hz!\Ի��^+��ĺ��� l�W���yZ4��ғ�ɸ�;M����C���ıCq�T�!�{ߢ�����PZ�(��S��1)��w-X2w.�y�Xf�@vX2͹v�?��E��e���~�y����R@y�B�_���=-m�M~�R�.-͞/���Ҩ�v��l�=��C��M�
��F�~��w����2����ik�F�p�N�\����=]��ϯSvka�ó�x?$���s"���4�NՀ�x�o� �x�
B����ٙ��v~��Fw���w���Gݛ�t���v��6H���h�S�����Sxy�k��.���)n�ʬGo
P�w�g���F��=ևv���ɐ܌�?wz���?�w��<�������1N���@��,3l����>|q����Q�א*E�}>U��'��u5���Q�����,�Di���BZ�m��N��"��|�m���]��1�Sչ"�M̘iuϊ�/��b�t�{���WvN~(�1v�5�~�1:���1��a�߶�"�6�KD�[���_���7�����ᡡ�l?O˛P�Kxf�g�,���ͯh�֍�]9��ѵS=�ӷ���<?�>"�_/��}"w�gs������G	�1��e�y*�v3��2U�*M������(3Ё���:�k6�_A��qت�?{^j��k<�&����t��񣤜�2����m�+������w�?��b{����Ps���R��B/�E5�P�y�t��n���(|��.��X=d�/�h�y핊k��F�����[&����r����'�7�Ϣӹ\�{ݘ�:\������n��,Jaq'��+�=�����Eݱ��s%�� �P_�\���8O<�ѯ2�F��1��R��O���V���3K>�8�՟�2X��k:-�,V�?ϻ��;�B�@E�ٕ��	>И���7��v��tb�(?�.Ȃ?O�<z�q��Z�[�{��e��^3���Hmۓ����B�ɆQ!d��X�܎*����҂ұ��F.aV���ԁ�M���5I�UN�-����_��Ɠ{���J�����j�T�gس���+������2�4j�<*?�{0)�����U=x��}���(�A�Th~-[�ԣ#��fȟ�%G��e�f��$�5j���]z�����#7:S�ə����C�A��M--�̳+���|�&+���9�e���/9 4/�ʋ�2=u��<`�@	��#��{3bc�E��;�Ԫ�(��,�5�k�Z�b�"�
���$!?5�o�Ϡg��Θ{�_ĩf��`S�Wla��-��_سk_=$�+����H��3ׯ�N�!2��D��B#��2�l���J��n�����mD �dYsn�[����J��h?oC%�튥db��K�l���X��+e^��'���\��%�oÖ��ι�����(������h�Iff�H����qt����|]�z���]Y�F�B�Z�ttƬkzN�����T�DԐ�&�b�s��<΁�bj:���fn6��;�q�,�7-qa,@S�	� ���h���_�ܻ�'cgcZ�͔ ���$�CC����JՎ,����\��`s���+�E	�̠��S�_�<(��w��w�6�^e?x~�9oj����1��ӑ���n��{������e�tB.2 ^_��!sU)�}�诡���K&��7w���i�o<6�nC��,Ce}���h��SC,r�ˑ�u������t�c��ݸ�W7�����K�{]�V���̊��܆���1������o�(#�iNp�};���ݶm�/��2�ZMfPZ�I�(� z��hV� 5�t���ANs���~:Z��p�c�6��,�@0�%$��X �����b��C��8��G�-�ؓ N�	^0@)�`&��c�e`&}Q���w��5��B��{y�)��tb�������AbJ�/���
?���{����?(C[4sfh�����b�pQU� �}C=f�u0��N��7�"�غ:��Š_s��鶈��S,��Y��O0�=�A�mP!�^�?�V%l�0������emp�7��I��k�>NL�I-6���E��y�/�t3�G��ƅ�������<�нzJ�`�3��ه�������5ۥ�O�-�#U���-��]�uˡ�#�� W6H����(E����I_FA����A����_0���I�o�=�|d\q�������K8��������_i�'��v��T�k�3<�(�x�j��1c��GG+���h�+Ԇ_���<��4Td𱋵>;ռZ̋��xN!�Ty�ק�c#ț�\�� �Ƥ���3p�2��f�����u��T��.[����Λ�)xEi��ذ�h����%ʮ��ɮ�i�'53"��9�p����af>15s^��-�A!�^PL|��1�-�lr	m�?�P�Y�`�6~���:���Rg�\}i�v�u����Z/b���k��Eif.f�
��8�T�xrn.�fWU26���ܗps����`��= �U!����QQC�r�§"����ٺB>���;�QiJu�[QF�z��h���)�ß���,^�*%�O+�����) �O����J-��A��(���#M���,y�/�tz��*:|`�1���nXY �5X�J��Q�C��X�A�������j��V�K^��5�A)����n/��>�l'���`��>�q����"���A�0�-C|@#�� xmGkV���#3~��x�laD�0�k�'����g����߲�8�'�+�D�|�>�r ������#r��.r�����nگ!(���e�@AD����_-b�^�q�0�����9
%B�*J)�롟�7��	5��F����CT&��u@��4��R!�|��������^~@y�B������K���G+<�R�\̬W�w�3#��I��r�.y_r��8����� �G�����M�fI�|\(���o��٨[',E���_�#����BCQ���/��[�Iwܜp.%�}zIaf.�ȍ�:ڗ5�ZZ@S�O>�@�}��|as��s5����ql�H/<������c��A��JZ�5X>ػet�I��kC�|����p�2�����Ș:o������D}G�;�����w-G�>�&�n��`tϯx�5���H��A��h���z^�q�?tv)�ǩVڜ��"�d��=���10
9�s,W2��ed�����W]��������0w^�C���;V�К����ށ��� ���嗽�j��H]�v��Į��8������p7s�E�P��+�I��7��ADlY�C�q�t�f5tb{q��of����/�N���8���|����"%:3b��0^k��?n"��>S������8.ZU�Q�6��}�4���'_q�f;X�R_IrB���f�����}��C�c+)��<G)��e�Tcq �Y����D��G���l8_�vO�?"���;!�d�|J����-mt�4�/oH���z��J�O���e�fed��������\Ǳ��mVtO��Ռ�� �ة�.���ug�49t������*a������LS8�
CXI�\߳����K3_�z?�,^Y�z��b� Qɺ�ow�]W���"��*U B�	��=;��SYI7m�_�i1��(��SV�����ru�*��x��<��zܺH;wlZ��?b3$����F�HT�x��H��\|1=���9|�B�y����ʱ#���:2{蟻�
����dG��G\�ܛe|�ɡ���f�U����G�iM��ӿ,��7 ����Om2��)���-�΢��V]���Q��<��������|*�8�`P��=u��gm�z��y~�@M�ibV�ֲ�'�K�B�g��C�\��:�q;p�4Z�j�E|f��s���"�C��i a@�d�.�N�C�Av�b�׾n�6�0O�ovz>*��&z���q����јO�Sx~�2�'��x~5��ג.jj]�(�fl���r���'/�}��ە�)�9_���D1�X)�$bn�p�+w���~̓
5�}7�H��_�-o©N�Ȧ�+��T���Rɺ*M��[b� yz.��+�/�≳��3�pjQ�����-���;]yEt�i��PIH�&�<yvȢT1���SN�j�rd�ĴT��o=74�}O���p.OK-]�*����j�Ë�B#<��-�$uǇ�]=-�(Y��4͵0���������+a�����2��q���r� �w����-��I�Nf�
(�M`�E#q"��#z�6���v��l���f�GA=�MY}rGl�?�P3_��|�t|�V���@��A>��K����Ҟ1�7�f֩� xɻ�>�'{	|���r�Kv"���w�<m)�.��y6cZ����~�(��$B_�7n�Ud'�7D�}Q�����%\,����<��7@�\��%i��(�Jſ5��Uj(�7p�]�����.��Ԕ�����#�ݙ����|s��Ł������s~~�lJ�F�E�ܵ
�H���3�6��s����IƫaL�"�ʷ�;�qFQܾ����r�s��|����y�T_���ޅa$b�����-�B;<�&��H��o33��Y���T�w��k��f��F��(���Ͳ�����f�H�G^ה��ͤ��G�+l|q��!*���`/�����B�c�Y��#"8���\'+�ޠYWU0�r�G�� mF䉘"<r=1Q_&3H��9�:�Z���ޜB�΋8�+>n�R�A�*��fRJ��ݦ;I �.��{�}6��2 �+U�^,k��Q y|�S���v��j��ޗ���"bѶ� �������E�A�kW��Ma���R!c=8��ef�~8 K*V+c���PC5s���?�����P�ͮ�'YA ]9�k̐'Ԓ(�u�M�b�\��C�@�+���6�t���%�-�N���C���K�]�gQ���͠� �����_+];�+1��҉B�(�C	��R08�M�K�N�+fN��2��8ϴ2O26�'�{~��vu
=�"!`�`#�5�П_ۜ�CW�C��z�}�-V�W��J�����Kr/��|T�Y���{trC���*a��p�l�-N��\!��"�A~~0O�h�Hxh����-H��aQ"F�hz�fVŃ+�/��0�Hr����̜��Fl���0@{2�dvTͭ�؛��|��n�.	!��u���::*ԭ�\�-�u���|R�T��%��vf�K��F�!!G�o>���cu�]�ё|�4 ��������A^���LLG-�0EB��EJ�;J�١vzn��t��˭?�6����t��r �]xZ�[��Cc������U�ÎS1��Uy5<Z���kG���� ������&�}	V�v	˾C0�[3��}C��r�q@��v����������Z{C��;����h�9}d������p|LVoѯKUKf��F�4U�"�SSNN.��d�� ��./�,�-v,�w0�`l>e(��_�Z}8�x��r������M���3GS�_m���6i��r��İ�=�+-�YCF)L}��/~�qK�Jјk��6C���_�eЕo��^|$�,�l���+S-�m�]��$yFZ>���T�S�az��'�;�b>G��R;h�pI�n��(���
2I�gwBQN(���8
@��N=T��j�Z�!\D'uV�% �cf��z���wV������cm}>~�[["�.�.q�����'$�n�tZ�q���\}����Y�v�ߧ�V�-��e@�nO��V�W=*��������l2Q�0z�ӂω��2I5}�`�v~q-���A+<?�)2)�3�w�H���8���Ȟ*ފ~F$���9�J��S����\���I�6����(_�便��@�Uh��M���h�E
��G앪�ԧ�4���թ	�����~l������=�iC}9Ġo�f���1��c-����#��i��mf	Z��S�.�j>���;e�՗h�m?���~�8�L�u��_��9�+�R>�]����g�Ƿ����v�o�dKK;��HA��2@��T�٥^�����H���˛����	����? �Pj�U��uS����,1��­��/MF�����@D��]qT�>1������ m�v@.rG.$U$f��K�0>����2E�щ���H�"Ƶ	}#�h~�2��iaN(lƇ���h�P�X[�Y��m��cajWHL���9�Y�tѻ2�z�ȅSY�6n6o�]�W���R�Nb�5����{5�^~}���V+��7CΝs�F��?�-*4�5���aL�׭� �����+�<&g���<��D��,�Kk�6��m��&Mo�0�$�_=�}	i��ك�*�^$֌/�TKn2In�Z�ڔ�lBj������M�����Vp�WB�za�O�����L\����ӌ_u�	Y��-����K���F'�M��"��3a�I�|m��[���|)��6,�1�X/��EsZl�>� ��}�GM[$��s,\a�ŎVΛG�-HN���X�֓���ID��Q�ۙ~�k����R=;S2Ѷ;>i�ҹ��c�� ��-DZ�Ng=��?�P���e�j��d����5s�^I�;@�mц�wG�Er̐�G0�����^��� ���5��T>�g�:r>���D`��lP9�^�Q?�Ro>�Lp 5Zf*+�|Y��7̘*��(�K���|.}Թc���� i���q���̗֊	��tdI#{��}p�������5��S�Ð�m�~����Y424Z��S��F��}����F�	ӿ�N�����Bf���th攟�{�"���ʄoU6�yZ�TXo��)c#$8"Yv��ɮ�W��f*j�*�~��ҽ]��B�ų��z�p�t*����>�I�%0W�uMz	N�+l���)�ێ���%�Jf��wՇ�3��3S����f�����J�C����\_��}��A���	��+}꙰�wGG���y�@DO8�0fP_(����t��N2V�0M�o���ޏ&��^Į�d^��f����Sd�#�o-�r�}�͠�L�$���Yha�]767_&9�,����P�.%�?'��M�H��p\�~������
��Hp
���>��{:��-c�x��s���i�6��ceD��gK���m��-��d@Dx��~���^=r���|���;x��^���B�@o���`��<��?$�ݿ�=�����<���*P��+�a,H�1�y�HVGn"�O.����}.���9fѥ�V��V�:^}'�"�����.T}a���;�Xw�͊
�k�T�4`�"���=�H��w3Z���?ɖ��s����.i����?!ð<����a�)�v�w�XT�~�[��S�c�0_}<����UԀ��ߖ���0)�R��>��l�B/Ԫ���E�IDhx�3��*�0p~��N�H����B�%�#M���+�_ ��tFo�Щre9��|���;zu>؉� ���>�;i����Lz�0�xo�̴��c�{�e��� �V�tNWG�W۵:c��ݿI�m�Kڣ�����;Ւ㲃�$9��䳦u�ן�RJ*kj��V��;������Zw�i�.D����U.iuO�d����J_��գ��쓡���bB5�u�D���N��1 +"B���2/���W��N!�4����H�t�����w���n�9�:>��_/��(_�& 8U�ER���ɦ�<8�=&��yg��2�������J�I|J@<�0���و��;l�j!թq>�^���t/i�^�/�u�҄5q��LAL�������U[�9I�ʁ��J���S�K�^�Է�b6�*̺�d��@E�c�$�AyeL��Z��Ӝm(�!"ĭ�Nߥ+�cW!}ݝ�o����(���{�t���l�F�t*8�� ���k4}���9V����ϵ�5@+c6��>�>�6X|�1�Ǝ�l1��_���U��uJ�^�x�=T������z�v:#���X�;7���l��+[�`�b��R yC��G-�+��Z�GE-���-�0!*��� '�֐���dw���xKs<40��\�}ЉA����l<�{���xk����ǥgH�^�}���*@�-a*���ۑi6ֽ��U�2#�`�5�Y5U�r�޼�/8J�=���9�2��C�W"_�2ҽ)��0�3&�� I _rՂ��b���=\D~FD�yG+ �Ug�ӳ��ϪU���R��=�[)7�˂�4���6�Q�u��x�>+3�������D㿯����s�����>��ꧨSK, ���b#�Pu1��O�'�E$ OQ����/ڬ1�T)����
pn/~�#A���f�6H��%U?����b��_q�u/��vS �T5J�.�=Y��k�f�*��2�����5�Dm�0ł���ҋ" 	M���&�$����H�z	�;QA�zBK(� $�v<������r]\"lf�^k�}�kf�l��Z� 5~�ϟ�_��jf	ٶZY�l�MX�8W��Q�&G,X�/[޽��#����c��>��	)\�#��_Z��/���a�y��Z�q�,�;Ce@��^r F����/���~&�g S�<	��"�"P>����d�I�`ֿɿ��Ss���Yb�)�f2)| G����w �����f�"g�P�`�����Kܟ�@\*t�"��s���Y:I��k`ɏ�B�e��Ao�& C�S���~u���4>�7�� -���JH?��.��~�ŹsWEN�d�:������W��3��6��X���^4ͤh�BM��ޅF���N2X/��l|�w����2���W�����k2W�"\�s*����k@��{A!��T�(��� EΖ�п�m��\�=_�1�@�iǆ$�w�G��~�G��Y8�p:�-�����Xu�%�ĳ��ٵ�]�~\��2I�74��v�d�)C~,���`Qh�;�c����к���|J�i9��V�v��A'I*ͬ	
���Ӻ���Z��f���nX�ȯ��~R}��rs�dM��WadU����z1p��.��X=�t _���恊�4�b���7���}��u����Pd��N�Y�TIǂN���Ӈ#���_��S��~��P����'4�>�cB�J=:ס��:�10S�^�֐N�'�h�|��)w�5��7��:�F>�MJ�ro=��Ϟ<y��k���3�⧁sV���RR���7����]O�`,� st����ؘ���͚���!�+O�Q���!����:�	��ʽ�k�"��;�w8r~�2��TCKi������K�V{$i���Ai�Ղi��bCR�WF�*��g���y=�t�9ȏ[�5W�@%���g#3v�e��gX��JZ�:Noz�Qۺ;�GĦ�A�i17Q'�fZ{������x�UU~�B>=��E޿�1X	����#��kP^��n�6,bV%6�����&}Iw�:L3&���S��6�/�~[�yce��
��x���մ�Y@�:�t�$x[d����D���܏y�����-~ՓW;��R�uu�����O~>%P������������ApN��})��ݻ"��L��6Y��J�eŧׄ��}ȹiF66��F\ښ�A5�L
������e�n>�~��-zMwM_n���L�����^����L	��eӇ�N�;c���c�U�HM��zrM�-ԯ��<�l�	��`d.�f��I��x�+ N8(�ٻ�B���鉛��ɕ0chk-`��!�3�W�'i��%/린+�4��Y!@\F�##�;�����Ȼ�л����i�a3/IR���'
��U����<!���
�����ˇ���\�E?��B��Wj��],|Wf߯ƀ�Mr0�^Ȑ�g����<_�I����=����ho�G�!��8�}�a��I���6��dv�����6+��%n(m�i4��Q0��셁�'ų3p}�$�	�a�$M�O�-51�����֬�Ϭ�����;�����!�2$:K���I�D[�@�Ԙ��dg��#�6К��$2�|��F|H��Զ��3�c�IuSK�*Г����
r6�]�v�6MC��P�+E�ZZ�ڕ�U��X��2�?��	�W4ϟ�#���l�R��"���l$���2�\\I�%���~3�q~'�y^�&.K�li7����a?�e�μg�mt�T����}�8,�y3đ����N�`r�{�9Z�ܕX��ٚ��{�(]'�6��cc
��ހ�X���<���}逗�_PLR�$����Em�h�&$�_���_[���N�x�(���#��e����5��b��1�q��v�ɸ��0��d2��O2-lZ�ar���N��Ӱx�bͥ�;���лƮF�ղ<�ۮ�dڍ"s��pM�����8��nYz{<�����'��gG0��[g�ߑ�*M��T����	����2M�=2䭜�KWe�O�R,�-�B0)��޽�M^��c�����$O>`w&��N���#�fi~S�z�uɳ�6_@ 2Q�
��^z�NN�OI������ۆ69B������J�W�I�U7�M�t��sYħ��0�ZS�$�y���e4Wgz�${�P�d�F��p>mL��J�z<����v.�d�:M<<�Y���r���H<B�}M����|Ӭt�=�䫙 �s�`��dO2��H��qF���dA)����XS�~������[~��[���6]k�j�ى.��W���%w�zN�?�]���,x�a*N���`�:E+��g@��Hm�a�n�c�@m��Q#�BRGA�g��-�{��������*�my����� ����g�̢��3(Ȼ$V��-���oF�L\�vš��/%�ڵg�����X�����j���\ 6�Զ&w���n:��s���w{6R`D$�{�V1�$��OW�!��\�����(��Vۯbǵ��c2������*�	��':P���CYp|vwvV�e̜�\�ϖbX����o{p=�DRrj?mE�X���Lyj��g��MW��ց\������wƧل�C\�R!Z 	�P#����w�[E��|�<�L�R���w��η��p��id����$ucm��9���'��-F�# /����8 �j�Tϣm��'.������m'0=Z]��L��霛~Ҹ���VF�������i�fF���UXM9����H:E'�-|����z���;b��"�� ^>5� L���^���NZ�wfƵ�.$iwK��z C�;�V�]��z`L��)b�g����@iV�Z��[Z�*O�"�v��F���W��}c��~����-�au�X	�
��������5X[ۺY�-���(:�����E=��n�^�a�恞��%Ӹ�l04	��My)�x�:�7H8��z�ae�UG�Xƅ�ꪒ'xy�O���<��r��o�HN^�1Z�៮a�M$6,��7o�H9BXd,ܧH}Zz&�7w�����M�'�-��OÇ�:��q!H�n�=��8.�0�P�	u:d�����^Ư������l_���g�� �Y N��m�|����� @[��W���3ʉ'�v��@]V���3�n��ΪF������Hݼ)9�2>[��<K�F�F�òa3t~=$�輓���z-5�䗗Z�-�����{/�v��UN� ��555iȹ�(�d���Th�MB��or�j���ڶ*����5�Ş/�0J6f��&u7���vC̊CI��9Y�(SG�^%��v�D�j��М���[���ɚg�[��J#QA�7��<KQ�0K�:u%~K�a^�����z�2Z~.�ڈ��3��7���Lh6S��[�B:���Ś>�2\��dS�"Fuj m@@Io���W���n����{#g�=[|��,�g����[T��L�[�F�@�V������;=�/���t����z|���ӗ]��l�½.Q�S�΁�C�j@�_����A�	N-�εüeH����:-1�%�Q�:�Xo�r���lEv��v�hg�3�q�}�īÌW zƛ�7k�՝T��m�R�RYL�z@�QЯ���9|�@���#o8��B�`y�i���#�ѦN��2M>�x�iV����H�ٛ�/�g�s8Z��MS|�*� &����5�|�5�Վ���g��N��(.٦Z�ͪz��V�����H�t����K�k[؎1C�E�����E9�-�˽��7���;j�pn����i��W����݋U����*�$�}
aΠG���ⰛN�$o	�:��O��Z�VI4�!WHur�	
ىߨ�[�R�3�fa�Q�6j�f '�Zi?�b=8��MC�Y>ŏ��*c����+�UX^�`���ۙ���|�]�rq�phǩWu�_Oe�e�i�88��L�٢�Z1V�'F\�1�Ŝ�Y\�C<��Y�"��(w��h:<x�pH��g�a�����CE�
�;!�?�f���j�1N�B��*��!h��?�}�x�
M0�b�o6�e0��g��żU�h!�L�`C�(1{pAw��ڝW�+��赆�IS���(,�Կ6�f9�רb�C���cԛ#;3GE)A�����^\~K��S��	5�~ �b��`�d����,>wvTw� ��NXm��[ �[�Ҩ:G �7v4CNA��DWEYU\s�ũ���d�����=�y�p��_��(���q
kU��;��m%N:�s�� ���EG2<�1��f�&��a<��fc�\�C�?/����H?dP-���G�h��!ѝ�ҿ]���w�.���ș]2���J��	r��1��&S�Y�A�pis=G)��.~�Jd��.�g7�b�砕tw�[zx��斒�rt�&&���L9���G��X"�O@�N;�\gR 턉S�̿��c?����ޣgc���3�P�@���=7%�
ٟ���z p�-��*�(�s��~���N� v���+�rR�r��j�k��8���ɩ�2�u��o�~I�+3��/^����)�F�;� ������6�����Gm��ko$<bt�5�L�iw"+�w��^���
���a$D:��j����^͍D��HӑL"�d4E|�bD� /�rK��Ǐn%�[]WۅO�db�#w����oCe��Dy�ظ�W�W�+�q �fy�s�rw�$�L'�u�W�vZ�D=��;�?l�<X��=G�fa�t����{YC�.u�B�����W�.U���q%jY�)�p�jX�?�-�{�״�����4|zؑR�Y�9�]Pr�8|�{}~���u+;��J���g~L�M�P\h�'���{K��L�o�Z���������uV�}�;*�����G'傖���AWQG�Z��4g*�['EDo`o�<n��CT��,��ol�m�^ ��������s%[,���9��_�;���&eQ�^�G�����������`ڲi&��6�냮vTtQ��>X��)����Ւ���� &��w�TM��8zϚ�׳l�����A6y����+ul�{��\�1�c�a�ۮ�c(Y7	{�׽%`,i�p#1Rn����ڮ�+c����,s�DY�GA�8;��_�*%6�3�]ܰ��F�w�������ڼ[)���E><V#E�tB�e��~CY�YB���#� ��LmXS���[G#[�y����/�T��u���R�A�e�a���_i�e�|�O�����b�NH�x�U��*5	�����I��K�s��J%s���ʖrT�魰��=�1>zr�œ�#֞�h,�Z2�r�e>ߚkh3^�E~Q���RJ|�먚����L(�����\�Ip$���R�o<fC���!e݅���<���"W�&��Q!��7y� �s�}��B�U���w��X�;�e�Da��f\[���M�cPv��X�~�;�U��.�I�c\״��4����1F�JͿ��h&�/��}/jpگ^o�r�ۃ���T��*��u��3��kREfS����W�/m*\ўyPZ�A:����v��f��Y�B�LŋUb���~�+T���q���w�ŽU��ݏ"�[)V"�4��_Y$f�|���So��/�+�����1��ёX	���M�������U ����������F��pG����|�t�La�=��izqA�h�M���G����@֫��s�vXά��*���G�Mh��٣s@��Kݎ�_����-�.f�b8s�V�a��qW���V��O�s� �ܲ�w��j����wgj�O D�c����u�[�&�Z�G������{���u*��0%Fw��S"�}���+�����Į0?�9˞R�YF�Fz�*�栖5rR�`�-�Ȯ����}�p�R4�RN�gO�_Y�"�
�d� ��޸�����׿ U�>���C�.+�I7B�.�����]�}�ԧ�VZLqF6�1D�1?Y�]
n垐 �5�l�֭ �6�jU͑��쎌����|G�;R�IBs�Wl'tj�u�yc\���v��RQX��I+I5�M����4/v>tLix����D5��j٘6�_r>'n9W/5���z%)&����.<q�ߖ�����P["���X%��w�2mn��.��wZ��\�Oo3���n��m���4ur)���8���������Y�c�'�����+��A�O.�%\A��AR�/m>*�L�TE�	�<�q$T�lo����npk~Lϴ*/�@�o֮�c�S r9��+.�4W����gN��&\�#*��!�����ݧχ�ʐ��t��VK��ϯ 	Fb�&W>gʸ�u1-GC���G��f5�P�['�#}ؚ  �nyy0�+�b�O%ҕ<��
�{z���c��0��?6�>H-�Tp>W�;�B{V���Mޮр�@i�}��Z�+A�=Sm9u��D�Nm����$�H��}�k��t@�r��{�ؐ���>5��P�$�:t�W�o���v�/�����+$�zc�h�_�+q��.����,٫;?��� g�+������Ҋ�T
]�t��f4+(�g��r;��ɝ�C�*8ݛ���@�n���ǣ�I�"=ml(癭��qb�4�?ؖj���%�}��}/�ne�9�2��5=UOd������Pw,
2jF A�\�=���|� |���;=��͐�b���<@�]E��d㒑2!����9�u��0�M�B~�ƻ��в}��p4c�9��n�&<��1�U��z�P�H��p��.t��3�ePi�*�������iQ&�\����#��E�b%��Z h�<^������y���U�=)�
�0�6�%�2�[�CT#��B~���w���2eF�qw�������jV���-�V�>�_������+����I�n�������v��?� �2�q)f5&.	���96tq�*g�;;������)�Ml�4b�	�9f��[]%�%���ID~?�%��e��8O}��`�]Az�3�3=�4;��������䒉���>��w��ѥ��x���eU��W#xÌNgI�Qr�ԣ�Uݵ�S�T K��'`�rEV �ɩW��d�����ƣ���p��	�X�(�5�g��jJ��>�϶gӇ�L8ow�,?��%����T��o�h7�OX��M�/��忚2�)��b�&>�����7�?��rE�쾯Y�t��z��L��P�>�L�;�fZ���<����c�#&I G?Y�!R��^)�b��N_�2]�ͧ:��L���p��=�=!��
���8�$��RD�as�ײ�#52���6D�}%ί�F�YHw��e{�l6����n�<v��X��A�'/�; ����%Q-���Č]I;��Y��G^Wa��Df����6iY�o�eXJП�-�a6�Э�'+��:�OAߪ�߬q*�k+�ݶ�uoO��gw�<]a�l�����-�'�V��ma��/�&��l��S��D���J ܎$����m�޷�{o�I�n�4d���M	n�j�Q�a�У�!��B����߻j/=$�UC_z�R�fuA���؝px@�fm�NwQ䷻ש*��0s.!#lɰ=����������V���T�ظ[q(Uc5��m�A7z�}�4 ?�ͼb813�ԭs��9 �G�)�@��C��0�O��p��~'��y_�S�)�&a5t�=a�ʒ��][�S�[Z(C ���e��y� '<��n�WTn��ǌX�����1�B o*f��-� �X� _W����d]X��y��I��]�6�ڎ�	�JNį&�л~&����\�oԛ�伵q�}oߐ5y��,��)�S-�;8� 5�b�T�5����|��8*݅��u�m�@$���t�CZڳ��L,C�E�+�?��C�3��s�5J�	�J�`��S! �+���_��*�{t"�Fg,�FgB�����%MM0,�U�˂+L��OP\�r�9�5F��듷�֓;�������z�ɣ�@	�V3��i�x^A��[uQI�/��C_��]X����IL�C�=j�Һ�^t�&9��=���<݄�?ߘj]s4�6�7M�9b����[RPh���+�k��Ս�U� �Wz��6՘*T+6�a�}"�}��6��O���Mk{�'~��'�m�/t�^Q���'!A':��_�!w[%�A#r���Bfͭ��x5�e���'��G��k��]�+��QH���lmo�ֲ�<�~�}��>IL%,Ư\�v�&������}3�W< ✴=��͙����v�3�����!H�����⡜� Uv�<O� ��o����T��	q��V6����6O�Kh��HR�L��P˖�Ϛ9Q�����{�M���K}�2�~�-�ʑ,�}�c�N!��\q�6�((\����{�:t�%}9������DW'9͉L�4�є.��d�؞��U�l���l����n?[���\����> �]�7�LiF�0��7a����}0��A�p�I�tw��Ŝx�Z;���Ʈw%-�W�/��t�/��Z��F[�xG�.����KA��֜��I��w�W'=�ƫ�<�s����Kn�mS���P��֥d��R��B(f�bx�մ����ﺔ�J-�0Ei�R±ء��ė>��)KB�XT4
� �6[��,6u�_����gb���LY]%���U�h�p�U}��=5>9��~��k��Š�j�ְ;�������_&9�-Ƽ�om��x���o2Aeգk�%��F����%9��a�緹���·��<��|�6i��ء����g�+�UV�j�O�i)&���y�Cd�`����ne�7�e�:�M�Yeh�Oj�Y�*��������?�q���㶾�Z:I@Fvz�r]W�L�����i�m2���ք�~�^�i�o��)u��,5Uw,N>�HՖQ�8�C��Hl��a�L�����pT��U�`�$��h7Դ�܍�14h��-�@�B(E�Gy�#יD�{�$3��W�}�����o���R��=)Y�l�=R,Ax=�����#
m����o���	{�W�5'�2x�c_q��O�bx��F��u��9wy��-��c�A
?G1T���=7 �~�A���e���_���$�f��L�2��]����f���j�-�&[�X�}>`+�Ԑiz[q�f�a�p���{�����RM�)�W���l@��|wP4ZC�=2B�!g��Z\<��gDV��=,��'~��K�]���m�n����/ƽ��*
���M���7�������
���n���`7���'�^���Јa�4�ı�+�2�ٓ��G��`��U	����@�9�n���-#ҍb_����x���{H p7�_n1���������f���G���m*4<37u̼;�f�t�jBv���=�p�<l�Wm{��K�u�z��1�|���y�<�a��h�k�t.���Cbs� /��Ԑ�͍��� _[�-*�!�ӧ<x6��q�Z<�R�������r��X�ʹzvC�QW�d�C4laYs�Riy�i^��:Gn�:�o�͕I����?�0Q%פ�x�B��ۢ��H���7�Ÿc�zXrSا�2t����A�ɢgn&����:{�,�m�+���U]���B>Wqi�����q�jNE)�ڈȩ���
4�I#��ٖ7(+�ي�>.!lf�kQuߘ�����L�6S�.���Il\W@ij}[ ��%� �<?���-��&�q�oɷ_�~�0���f-x�ں��;>jc�\�X���x�vMǽ	Xtk+��0���t�.#���?"�J�{�R��D_A�x����f��n��5��5�=%@�'�!6`�0#[ ����%�����g�#S��4���(+�S�G�85����G�{��Ù=���ܠ�09�Q��<D�n�=��0ټA�|R�_x��-��,�NSC���e3S���U.�R��!%���/�6V����L�з/��Qm��#_t��u����TM�<�8�
���Q���=<�̝Ҧ��@D���3$��voəa�\�ٺ�����ʙ����`"l 聛���e��S7�* Db������*��azn���h������p�iL��'���Bۓݐv�g�5�^�>�W�F�,3㻠�:�!���$F�xL�&v�	 vZ^0 �U��.�ʁ�"�wp���}�Ԙz!�H;G%��4���Ia��ڍm��[��K���-�w+�P���v����6G솢�H�}#�=����@!�V���)��L�?��ۧ������%RyCi��l�9f�Ӻ��)��pg����J�Cxd>�ܗU�����(���CX��JRGϧps��"��~�7�5ɻq��{�|�)�B�c+-�MP���z�a
l��/A}�V�{8k#��
Ȓb���k�jn�Z������p�k�Ej%=���nPB��-����S�,�\]��Cc)m/<��,j�m�?�{z.�� ¬\�6���D0k�f6�#6�~��}6Rg-,犗7����-�{-;ɏ��-(l4��p�t o���}(I*4�,�4\���]��Q�a��HXn��V��
��~�g(H���E�U�b6�\�_�6i��-�e�`���)/msw��Mڔ���&݄t�W�����l�� +���)�
Ц!��Y[���S�U���_�r"�����b�|#/U�ׁ5����5>z�ю��4}��k����[���y��v��LC����k1V���[-�@�1ٛ����t����gm~dm�n��Š�aT��E?�j����������C��3���� �k�ʲ֭$�Jz�W���.���Ϳ�`<c�X��|&��|�G3�*R��7�6y{�?P�2_z6uu.M�j��u�n��fB����t���v��;\�17؟f^�Ì�~u�����3���7�J��m��w�����ZS���0��Ǧ�lK����R_
���"��y�Ց�:$���c�p���琇㐰 �K@0���-)^e�N�׋��%��Y|�a�K..I�P3�rK��.�a��V�S	)gЪ�ɓ��4�3��Bu�[�h�vl��i))��T��!�
��eXO�z��ND��Q��k��`�5��{`�l	L��w�B���\l���5y�v!w�e$Ow�Q<v3���hˢA2ܫ#n��\�2��N��l�{�'������w�I�/�0�P��a[�̋Y��.x�Ůi"e
?;�}�ȓ?���\Cr�r��i[�R����e�p��=�:e@��;�F�B�Z�8m�,sI�QG�b����}��*�p�W���I���Є��B�6�'���a����'o���d>������(<���FC]�㥥]{۔<$��K*�v�Y$���'�3"�e����X�#x,_~T�f8���eGGF
�K��;<��&��J4�&�J�Q�? ��?����=�̻)��]k�^�$�O�4���y�b������;jP��a�%��� ��y�>ީܒ�%%V<��p��<�xx!�,�@6I��>�Tǆz��&�������:���&��j���>���8���n��~�������+�<f/����-�����æ���x���G����pEUE���#�9 ]]>6��ld�"u��0��H�J�B��H]�᩺cA�����,y�M�	B�Y�A���RA�n�q4�`i��,�C�����n�tlM�&�`��rgT�8��y��i�ت�H���kl���Sf��Q {.h_ʝ���[C47Y��J����X���$�Z{q��ᚽߘ�<wgY��z3�(o%!�����������m��z~�t�)�@:��e����p�C��K�:�3��H�����e�umg��t�2�o�|������`�v�B�3z����]d��i����+����JuZ�	�A��4����&8���/��@U�{��D���Rx\k���*����-�<%�������j�,+�<���({s�j��k�ιm�6�ć;�5��X`�����B9�)�ŝ��2����7b��c��D�N��=]��#z�9Vs��cҦ2bq�q���ό�B��
�ޞ "n����:�h�^�8��-���;��
��Բ�~�HW�6����Dj�9'�&�YW�.��U�Ȥ�!�I�'��C�8	Ɛ�ކo{b�5h�Ì}�jB�,~�%$k�C����B� I�ձ�vH\�5'�e�W3�G�K�g�����~�>(�������L~w��aI�v��6�t�n�CB��-%��)K!�Z3	^��i����%�� ��-�QK�8i�;��1=oō��M"�{��g_&L���-c	�KF����U[!А{���կU5k��?}Gך�Ҕ䁒pf�ھg�8�i�����W�j�f�s�[���Сx((3	Gj�g�e�=5&�X��n���.��0�2�ߖj�47/C6�:��
�@5^���۬]�
�vҟ�۟��~Jb GB�S�g�|83ks����
Z+�����0Zn���u&ѥΫ΃|#B���w���t�k�����D��.���^�������s�[?@�^g�~�9ݩ��̨VE"�m�
5<=��`�h(�@t������g:MAq}��tf��n/�=��Н�YB��*=!� T�<�;�.�0��#!'��!����n�,�D������&���jȠ£'�4�i�IK-����zD��dmH�2F������>�c�ı=M�y�	�76�-�a����њ.������y��^�*7N�a�T�f�߫|�*�IC�"��Ul���7c՝ԦS��E#���Ke�
K.���]r�pK0{)G],�ŝq�!���G��~�ք7]k0 �P�ʗh����-��)b`0v�G�MY��}�,��>A,@��� �1	��8+��w���V�U���Et�5���/TkK`%X�"��]��hh՝�z,�1fX�����O.��H�ӓ-��;�G�t��f�o�t��e/¤8����r�Ҭ�.����UrS��4WwS��|��[&ێ�0��u:��yNH�釺�&���OW�5	\�������=��/�^�^0>�v��2�PHx�7��o[ո��ppY��╅��_U�������GE)�͌�\n�t�D(�1	fצ	o��RL���ә���1��o���C񉆟�l����GR�E��Pc��Q�Ҿ���dйt�0���C��>(�������b�DxxTt�*���}��n=�]49�Z-hnDޯ��c4[�k| �:��HRݝ�$E���6L��M3��m��m��X2�t�J|�j�z��'��*�n|����IL;D��_���0[��0z)�,�9鎈|
�G���x:�3X��Q�a�B���1����~�-��m���1�'��y�{$� d���uT-��f�g4*�='C>�ͺ5sI+��l�Сǌ�z#��}��rl7��"�l/o��|�� ���tK6���};�2@[�y��'�>Pz�1��z�|Z��OkZ9�!w-�@�t�N�R�/U������z`�Z�����l@d�
���#R�����C7 �t����G�����w�W�uɠ/|��e��7�Vrn��!*v�+���r�G��N�9

�#%7���F:�g$ 1�J��J]!IR��灋n��l��v��4�R��)��J�m��r������U�e����6S�9�((�]8+�q������� �eJ�@^��I�����ŠD�f�#�KB��I�p=�;����U�P�<�&`T�V д���.e��yv�����k��� ~���;��i����uSɵΘ7?O��*�JY���qQQ*���B,��z���6Ľ��\۱-"~I�,��������ݽ6�/�0t�Г?�2�gm������Π4��4��ߜ|�;�ݬ�����H�m�^ mz�1V��p�#�V�f��6�τI��:Qjb�5x�����2T�I)Jd�qɐ|�zw�\���"�R$�V��hK�8!w+N�(��]��U�����P�K�s��X
�1Ρ����w�?�}ˣ/���.�zrI��d�U@�O��{k��6*D�ͪ5�պ�B���qtpD��l�@��{�6�z���T��ya? Iy7���>���ϊ�3���l��r�Nbz+�	4éT6��L���RP�
O����Ҭ��
i�"C{���(6���Ŝ
J����єCJ�k�nq��޹i�.�p�B��:�J'�P�w�>���+�ses��˂M��?�T���u�^_Y}WOP\>q��'�H���iA��ܨ�&����o.S�?<�@�+�Ҳ��ɀ���h�m5)���SG4��[���B�o�;Q��p�.�i�!;�KԱ8~��_^I�g�������_<Hv�� � ���f�?��|hBh̜EiFY|c�;����)�J	 �������U�.U��J+hUM�햙^^F���Y�7ިa�4&�$JS��p�-�УUOP<{��hP�Z��1��s�#ot���"�͕��AT o\=��]�ס븏�l@����0��^�O�)��"���A=�5�E|t\�\�J��V�w ����x�Q��:�Fe(��Ĕ�������w�~�;6)"84D�����fV~�r�Vde0iZ� �)�u���[Ɖ� =�')>zJ>'����4a��ߌ��ޙ��v�Xd~D|��Y���R���Bb�3���W������6�*hS�U� �R��s�W�Ѫ9��31Y��!��R��8��`]��kh�A�����p��0�%{�mh9���w��~��C�yRNP�!�*:��xl�x�Rq��'�V���ct�®~������FAX��R3">�tg~J�4jR:X��dC�;#�q�Q7�ˏd��7�~�6�c��=�6r��dK�ٻ&�_�����J�o]/��Y*��F�;��}P.�dq��XТr��m�F���l�Ú˒=!i��@�[~bN�-HA���]b���턬b�s�:�"!H<5��ϝ�����:HuU�w�mz�V�S�YնS7�m���8`��X��:[t�Y���$��ܾ��X:w^y���ȝ����ڈ��M��3�R��e��r��8�r�P���(�|����V(��)�>�j�յ3qO(KG��9�=`9U���n���&��rJ�R�]|b6�(���3�]�q��ԫ�J����l@S"����Z4A�Ŗ��}:C!{����Vn�z�C�ug`N�)F3�_K�Y�k�R�G��L�U<JQi�z�,�n!zB�O_l��H�eht�;yCy�ƟH��^o]���p[v�vn��%�cƳ�7pE�_E�C��SuL���_�Z4�=�y��Y|2���Ƚ{�9K���_�u�9��+�t�+���	��~g��'Vȭ��c���\F� ��֔D���f`�1d�,��r~�$	Q$��ц8���{�A��vq��uW�J^�Ec����7�e4�
۱��T"���ʧ�xm����-m*5r�(X���ǯ�=�	�N���~�U|����9���>}��R�d��R33J�u��]��W�YI�G�vd3$+�*o�S���|J�\K���cv�:�:5(�Z׿��]0�l��,�<湥�Ņ�P�G����<J�� Z>W�rK�d��1�7����!*g@������Cƻ�3t�F�G���o�;թ �I@�یh�'�)��_)"�U|
,��H����[*���X5��>��9q
�8hR[;���tF"{�;6���p��������qW���Ñ�'�Z�b"�dz'�ߣ��R�zJ�n��Z��2]�8+p�-�ǻw���ƌ��a~��~���ҍƲzV1V�n~J��9�	��yz��{��Z�cM0>|X{����6��ϯx�W�8Aj�{2Ua���S���Pb�y�@W��/�a�Q�p#n`�p.��te����vtvN(���9���;�U���΃ס���)��xZ�8y<aC��r����lm�b��s'������6O�&�;�V2�2�K����|~�z6��>R�gV�%vb Gq�����0�={�Ǖ"S���SYU]!,ˉy��� c���u�=u�e�R3x=�zu�I,,���xhM�gT ��QT��z��g��m �:wܛj�m>ٛw)W�� Y^���9�o@�cV*.��D�|�M�A	���2ԁ�ɺ{��W��Mlc�To�Wa��g�$�.�;����<�I����dke���|Lull�?J��i�s��h>�w�'#�c��8��V���m���g���8�����Z^M��Y��PK   ��XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   ��Xx�آ  �  /   images/0fa89018-bbd7-413a-af56-bcf37033748d.png�b�PNG

   IHDR   d   V   9P3�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  *IDATx��wl]Փ���ı��;�$!�З]B�e�!!�Z����X[ �(��Xjh�z
B'���q���W�|�y��ׅ��1�1ҳ���sϙ�9sf�;v�"r��Q4����OB��d2�A�pX��������Beee2h� �SPm�w����AZc1�F���lw���gͯ���'���J�$��СC���(�
����V����ѣGk�A5~O���M���� (�LJM]�̛T!w���ژD�!�%c��@�Yc' D�� &���J̡�f�$�J� 9�dڴi���k�HH�%�ɖ�[�8��cm2gB�������&�ׅ_Jk"������"��ƍS��ر#�x@����,---����Q�F����s��(�����e��s�g�J���=%�+��t�F#2n�U������TW׼��9眣���#�t������Ν;{Q�,���q����G���D'���J<��3��#O��\j��U��D2%sgM�yN�x�6�.�U{�HA}}�^�1j
p`=z����D��;}oj���


��2~C:<�@<�:oy<nj�r�D�FP'���xO)�J��c����Y�ُ���&�]�k���R9�/GHqa�4��p�;���TR��OQ��E\���㠃�M�6�y��db��0����WF���K
0t�gȤI�䭷ޒ�7�9� ^�l��^�Z+�s0,X X�����k�Icc�^�a��)S�s ��ɓe׮]
8����u��R��dZ��=E�>x������a\�;��΄�̊�
�6u�v�����}Q����v�y��d��@�nDR�N���uee�2��?Vi��_}��Jٺu�Ԍf����/�k��ʅ� �3�pHݬY��.����z�lu�m��#�Pp~��'-Ù�Z�/���V\II�����$۷oW��~����'� ��:�$262��$[��#�.�<�={�����|��r�7t� ��Y)����ŲaÆ�
���R�IW��t�I�xE/��dƌZ��ŋ�ꫯ�-[��ȑ#�1��\s�5RWW��P������'���=��	8�Ct,0$g���*Uo���p�M7i����ɦcЙ�������>�ߍ���rX�H�����t\J�c�jk��Eb)�u�2z�8�YWf.������혅
�1��=���Çk/E�ظ�� 'NTFқ� ���3g�|��Za: ���)�zP*ꩧ�R�2�Db�>$�:�l����7o��"�^�����UR�����${�w�R[�*��������:�*<q��)�g���u;!��
�� ��3OQ/=���F��7�Ș1c��W_�?�P�����2w�\�Ρ?C>�`w  ����`���OhYH��T!MH�������߫� ��~���By��������˵��N�!�0�Fh������Q��'�DNB���)�؛9`��i�����ʤ�$�7���8Go��w�;ϢWb��a���8Gg���Yc<�c�1Á�%v���y���`?�f��A�w�|�f BŹ���7d�Y�@���{~y���ٝO~�y��=6����<�v�>�����5��@��h��V@  	��_Ȍ�}A�f*��eo��s�.�R�jh���3H���3�����[�N�*}��eȐ!q�4;F���a�t ���V�\�7����}���g��=;���k�������:��h�B�vn�����+������[Z�=R__�.-�N*��V7� ��_��{���l����F$�V+�9{��1&ӆ%��NbZ��y�%��__y�7�<`�� ���%�tx��kd����l�j
���I��y���-Z$�����X��D�K;�Ԙ#,]�TMG?n���@WY�.Ԯ�T�I���D�MGr��v7��<��꒒7�ٙ�PnA
p��1����u�D
��!��A�U_A����R�n�]��1
~���β�����N�@�F��p] �@WYQ�����đ��`��t}KB�w�J�mj�ۼ1[�B� �HI�jEX����z($�_���Z�}�a��ݚ�N!��ȧN��0s��1�L-��"�8�c���F�g�H�z �b<�p�MB��T;�t]�S�O�&�h�/��!�U�x�͍2���nc�t�j�J G'>�^�p�_�h�E�Ĺ3����Pi����(H���� ��d�S[AҰa�tn���q`����7��$!X�
'����g��'(�8%�*D��2p1+ʎ�h7A7�����J� ���O���O�s�N���z?�p'O�&9 R�jjk%�L8@
<E�^���$��MH���<����('��]x�r�w����JDM�t2�-X%' ĩDʣr�<����C���̘��vQ��Ia�С2u�Җ��o�%Mn��he8˪f{��@v�q>�cQ��I����!�|��w���W�X�Ki���.;d��p�PT}�P�E�wV��hHvn����~��<@��K.�D���kM�Aך�M�4��[^���[/���7��u�� ��]�s�YH�2��866�&L`�-�~ވ��:XY�l�dvr�s�@�$/��� �L<��e޼y��s��k)@�t�JD�ɪU�T@�}��&Lp=9_d���ى?��C�p0�$�ś�ER��x����#���tR�Ȕ��$�F���_�e>q` =F�YZ���<�TS*(K�,Q��>�leL!���3���` �H"��aB�O?�t�T R�,^��'�����娣��[n�Eˆ1䈑f�`�j!��I�ç�=�#%�c�~��3I��)^d�& �St'Y �"�o��0��=��)���=�\+GC��d<,lx�Vo��F���p�u��Ҋ�l�>��-S{��,�@���=CR�)0lĈ
,���V�0Yɠ!��z�6!�Z�%�����i$��y��B	E���"Ub�$�~��",�i�q\w饗�5�>I���䈑� ����$�����2��"�{  ��%#��9 �^$pPa��zc|��E}��Hׇ� �6n�$U;wHA8�ͺ�C�a0fӀ�{L�ӋmP �#1X3�ڀ�`^�/pY̜9SA`|���A�x.y^�w��u�Yr��kO��$/��b��{r���"��ޛ��Tz������ԛh�������E*S�2�"�Xs�3��'[^`A1�[Ќ���<]3ۿ��\/4����몺8O�Rb�����{UK 	 �9��*�sy�<#0zR�0�,4����ď�q\3a�SS)7!\�a��V"����eb�QYݨ�C���H����-���7"�0��PU��ެKT��٨],D �Ct;�H	����]W�}����M;�%��,���w��x�$Ԥͳ�UY�
p�H�!�[��Te�G!r��K&M�[��1z%!h�X<%�u���U7˟�gd���I���L�Bɔ<��/r����������ĤPJ���x �D C K��/~�Ie��as�\��W2��݊�Т�X<-����'����	�L�������+�5� �e�[�~�i�Rb��4az�Ԩa4��%ݭ�#D���L�2�j�?���GL.�3h�\:�*7��Q�*O~�NVn��1�C�Y��Glk���sp���������"�gT�ۛI%�i��2��^�"���rihIt��u���
�	���K�p�l7�_Is
��< H@B�	�J��ZJ���a��R��ܴ�(����c���=A��庽ݚ��x�9�sލ
�vi�5�텲���e�#%���'���0�`�m��{� p-�;ʲ}Q8G�|A1<��%����En�G�m��M���Z���~+����*q<)T�E:�x��u�����&HÒd�`=�5w �R }��u�2�� �o�@��܉'��Q��>�(�,�qm�> z��գj���ϒ	Σj���[��Z������ќ��GW~�˭��¹��L��A�2~�89z�Q���)���U�P(� ���\znWAz9q��֐���������ō� ��}��-NnLc&�}��w"t�G��K��id��1u���J��z▧cQ�	Rτ�P"��&���m��M�A��fI4g]��4y�	�:c�\����D+���Sϧ-[&�@����o@R� ���bׄLa �T��QI�x΄	t��T��~K`$�i ,�v� �����7߬ϥ ��$�D'�#P6φ���'�LK�̡2�x�;
���Qai���&����e�kO�NH��X(�z�� ������0�Wr���M��q?L<��<����%u�DٲG����!e0U��[il�� D։�j� �A"��`��ak�Xs���C��:H����,�8���F��7^��~�@��ր)����S����VC�@���[IH�t,�ض�@��'0����q �L��H	�[m �<��Q��'�z�\�h�m�a1v�D�%����8LjQ�n@{eo���霅I=������0ö����%�E"x�1a���r�e.gۆ�� �9�������~-�5�Ȳ� �&��vl�.���ݮ��裏�s�����W�Q��5`���{�����*b�~���1�����U=�2I�*�/7VuU6[�;��wk��R��������/>\"Sg�|�>vr`pF� -|�=���׸ep���v�m��Ʋ|� z�G�3_@uuLHd&|&��;ԭ�Z+������Z��0T��&��C9	aK���@�����xUF]�A�F`)inK���$�e�W�t�>s�`��'��A�i��E)�!m	�on�+[k(+�,�����̲�q��iji�������VI���-�Av����xf�����	e�dP��($� %DCa�<�Lj��6��D ���L�QW�.(&�~�r1�fϑ��BI�v��?�\%/}�IZڒ�#$�[��ѕ�x6���/|��Z�~�1����	��:3	�mn�D�ͻo'@pC�+΅�'��qeY?V8��b ��_�k�,[]3�7���kss�C~#4��X�~�㨓���oм洙������QS$R迫�� L��$�	��ф10.��F=Y�5a̳�>{5��Fi�Z��S�5�"�).w]p/^���pvi�@�9�3���x��'3t~[�pa�v��|�����w�G���_;�[kiy������Q��͒=�X������J���H��uQ"�񑁵go  `�$�n� ��ez���Q�|��ڵ�X_���?����i�rfN�[�!\�^t�Er뭷��%K�] �r�H&�ʮU���]""���j,�"���DVo�r�-����8�1��^#}�Q�%��8��$�X#���HVV0�B�f��z�v����%8KC�#�m\o	3�I5��Ww˨;d��Z�xp�n��[k0��6�[b������N�l��i�{��UW]��I"v`���n[k[f���{l�l�+ȼ�6�z���.���R��w��֨{CΖ� �J��!٬E�M �8�d��K�gk�MfI�0g0�;I�az^��?^N��1��%'�]��T r�P��00H�`5.D�-�X�3�r�0v�����"�$rP&�����I=�Y�ڣ�䘵����`N��e-8L$]���e[kpL��Z4�2a.�d�W&�0�,��~+�]B���=�\U+��}ѢEz��|�J�'xS9��=�7+,y@��z�ˍ����>��蝌aD-	�K �t�Ac|�X&]�!0]��G$�����L �r���Z�`
dY3�}�˹�Q�0��  ���]v��C֤�e��m��� �; .�!�R�����O"}��i8/�B%�Q���@��T9]ԕ��|GO���y13�M=�v03��U���uF���\y�
<�E���^��B����I����6y�����z�+���s�D����}		���#T��l�&1�R��n2�KQE�90�K�]|�: �r��T�] G��LHΓy�]w�u�'���@:� ��x��j���8t�5�l�`�kj���4�TE���-��=��Z#��V6&�����/Si�z7��7�y��ζ���ߋ�=���Զy��<������:���s�z�Gԭ���*\k�e��Rq�iK��k����(;�#���K&��sly��[*\y�|��ְ}sm֜�d�/�4g��z�s~d�#) �����%߭5B�l"rMcL��R#����m�M��=���"ok�T?���9(�m� ldC��M�{E������l�o*-�+�� �DY÷j[�<�|���~d��R:�2[(��`����2z:�C�ڒ�j���&�g�o��愺��X.L������՚�$SU��(2`���P�O�-������:ɦ=>�d��e�Y�b�T�5��w����%&c�wy�/�C�C`��ҹ f������d�j�3߹�!�B�j�Z�"��l�$�2���zў� ��&���0im�� ��]e�1{7���{�<��2�ii    IEND�B`�PK   ��X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   ��X��MY��  �  /   images/6e704699-d8e8-4ba8-9ba1-d4b639f353b6.pngtzUT]�n �`	�ww�����mp��n	Npww��apܹ���xzu��^{�쒯���P ��O�>��H�+���qm"�}��Q	���!:Hk:��#����$&���GF\�0�4ޛ`��P�~/�������B4�I`�&������n��]�9"� 6�E�|ڑ
���
Ǹl��:�$�5e�m4���>7^?�9vJ�_��a?[�BCCv�!Dٲ�"s���#�6�Ķ� �5��Q��ߙ�0�o/lF߶�&�V�PP�<lxk�ylO,����i� =�0�#�!��yU���T��gBy�zΐ�
�X�N��]�#h3�5�\�񶼷�b�l��`��� ��
���v��r�Yՠ�#���O�S�L���!�i�%f�6sB���y} >�Xǔ��C^�e̜�۹e�R[��8��bT3����4(�V���������WId�RPɒ����%�* Yr:k���H��`�A2�N_�8i��/�9��J���#dI���%.�~�bA�t��B%�/!7f���q�!(�/���Y�ǥ�"��p8=5=�*5u�ʠ�2��q�$g� �� E�Y%��2�L��8G`�$�:[Q���NP��E@(d'߂�wr��#��WDhP_ͰMܸ�B�>`b
3�WnB�_�?�3��&�����E6�N�7af�,^B�"��f�W��&w���$�F�L�[z�����YJ�;]�k� �9,A,Ta`�F�ot�i�m{_ȟј���(�?�ͅ�^˷mYa�t����b�9<:-"���G4�%h]�($D	�hoB&�������/'����3�?��ޚbI��6��;���1 D�$�r@,���r���c$~�30\���$���C��8�X�p�i��u3hK
9�;�e4�Y��)�<�����_ ���;�w4}�����2�q#�4�$j��7�՗���}�bK�}�p��}ZX���/F�fJD����Yg�g;�r)8>MȜ�B9=?48�����v�
�)��V�9��߽_����C�׫� ��e���Nû]���K�S�i�D.��9�߹w.D��3�1�u�,�GS6I�6�ڪ�1��z���2+?d.X)�+�'S�	N��M�"��ú�_)+?��w���IEP�5`���-zM�BQ��jl�#�Hf�\!�|}ڲ�:�藀%]�D¯@M�(��i!Ĺ��U���:�:���U���L����Q����XI���ղ�����s��!���Z�9��wܷ�[\tTu
&>\�W0���,��QP��s��L���^�;"y�3����O8�3��������j;o&7��jw�R8M��%�d2���F
]�Oe&n� ګ��C��]&ڐ���&�NrCg�`}Xy�X�&��#��9�/��j�Rc�v1�����!�?/���ک�����͖��^g���~ѣ���~hm��^/��t'Z<i�ef�y�ˊ%�����)�dlK��)F���d:��q)�?�'ݿ\�\�Gon�dba0�$wyݢzW�{(��G4��d(���=d�'��ɜBcebB���Yju���LY��s�4ڮ���N
3O�2�ے��w�Fܟg����J�¸�I�4o��H�+��u���9_5M��`�L+�j���7�"`�������w��蓻�lT��iJ��h��Q�vaP/,9Α�Dq�:���YI�v��ƨۭ��;/X�+�}^|�c�9��L\c}�;c6�hh�^O�Y=�Lh�G��Hx���a)�����{p���:6Kݏ�/���5���e�Vc7��|;ܸ{��k�ϞN���7iA�!+�[I�؍�o0�Ũ�ϖ����4^�\45 �cS	�@�F��uf��>Ve��j��D�Z�>h���r��:����&����/ʍ����8���g��۞���3\5��u'<�aG��r��5�IV���(�Q{�+\<M���ׯ_-ll���^!�Xr�/�רk��9�O�_�S�#R�˿:������n���EY����4)|��K���i��bs����6�|�y��5�m�x6���÷ۏu�J5O���_?�J`5dƨ/��1�D�ғ��|�#R4<��E�~�F�LJ�P�����B�}ك}��.�K,Q��	P.�|9v|>k�M
���NrEڶ?mq�1o��m�=/��s�i}q�Ѕ�?����!\�(�Ps
�@�iQ:4IP�������Z�-
���XkAX�k�|�K��Y��o�je��ݿ�g��
gꈾ�}o�����23�����zf�IqJ��/��ֿ��B���z8o0M���oV^i�G�6�"!I�S���g����P��#����hr�����Ϻ���ꂏ�yD���p|cf�˹�s�P(w���!�c]&o!yB���.�}�w��E���F�|^e+�-g2½���c����
Q9�rx�ta4r^�}��� �m�Ԕ������P<y����P|�-''�)���z�K���|��'��6��,9��p�X�wS�UgkZ}����^A��RW�����Ѯ���*�ܞ;�:�0�A6�P���6_/w"�N���ҍ�2}��W��yyw�x����8-���鯚1�È6+sPY%���/x�ץZ��Oz��q#�!0N!�F5�F��_�Q��Q��(�8J��q-4mH�	Sl�;9��X�D�j�5�c-d�䵷g�� !������98���G���bOSш��01��9�=@�[Go��\���@���1eKQ�����i����{ �'��7ѽ��_tb����+��y��iI��Y8����ţ�uژ	h�@�[�aD�	0Zc�r�f�m��a)�x&Ӱ��gt��P[( ���˙��É��D=�A:�h�����K��u�,���Ӻ���u_yzz��mB����lQ���|�+`���5{����TLP[' -[w���ޭ8t$&_sɕ��Π�_�]�gQ����͹܀��C<��F����J�B��c�*����c�?����b3BC�zRنʦ9�{u�\���Z�V�+x��a��+dDf��ᕨn6|;�J{,8=f8,r�4Et֕��;ܽ���Rę�C:8�-b,�8Wf�Ջ��$#�&s��v-�9�R��	 Kw����j�>̔�S,�,5�6{(�P�(�\�Xz��GL��@�?��Zk�7�<4<l�:��������������T����h��1&�|�EWwx<�*���1}w�N}�������m����
y
�����ު�ΰڪ�Ӹ�PU��h
SRv�(�}�N83A�]"���J�誛����i���b�����zzz:����^�~h�#�>�6�P�G���)*��J7f�O�����Q���>8V�|�:�h#���m#�ئ�����Q�l���Jcc;�)g��G\��E���͏�Z�z҈�潶�b{�p�0��W� �<�'������dE6�oq>����/�TH���FN]��R�X$�����&8�	k�[���;[�8���K��~hcͦ�0cy7GhN}�,Z���j��8�ٷ�����㐴�.h/�B��L�]��%(:���_r��1�񀗗*��0��S=���z�]�7�0��İ5翤Z\Z/lI&��{0��#LFZ;�#J֦�V�Y-�Jv�55Gb�3����n�>�϶v�g65��
�J( �ê��	��XO�Ozj�^�klLA|���:�^�� �b��ϑO������>��v� j��q�?�n�"��e���X�8��0�/��V˱��� �Hg�����^q/��ڃ!��� ������[�Ewb{A_�aGd�p�J̑�2?T!�w� I�+�nB-))��>39�g������a��ni�2]�k!���$א�P�8�F�Q/u��N[K��X�=�hd�ܤ=��������e���D�o�.�.\	�{�L7$fjT�%��Bُ�M-��JrT����j�/(��4W��M�U�sD|�o��8�n\i2�F&����3�ug5b��̲�;#1�~��=W�a�;;���T���cu��3��S�d�܀�6Å}�I�x���м.Kh��:�6.
�N��>�#!<�u\Hbd�ٙ٢�𣅄����`M�'}غnޟkd:ct[8l�Fc��q�^tc��Ew.����ģ������k��t�Ce5F�d��y|T~~����B����CN{Y�h�1�P�2�+z,��	L1~�>zR�����;��3u:��7��/�eU�5�s�c��FK�e����ǒ"�ݍ�[��f��H�}��jC��[-�^�T�d��j�}���*�b��2�k-�����-zs��R,1w>�Y_U�ͤ��d�4��ܔ�f-J4�B]KW�����Ա6f��>���ze�<��������aK�d��l�㊶Ɍa�{s6Y͹�]&�$���2O��P��}5L--��I����>�-��n޻�IR��=�h��][�����d�����b�h5�԰���|4mgm%G�Vh��C%�MЃ�x�J�	P�#f�Xy����4�B��Ҏ��RU�P�����~���YK����k�e0�M��A��yq`ۯ����3\��]�v��ҦqX�����Y,���D�OdB�9��9V~
��DC�J�~͠��Nf�Hň�E:��[��b<�[�L�I��B+��S�%I�S�]ed(��c��+V`D䖏N��$퍦�w���$2�͊��5~ŪϮ-@����i�T��@��`<�X�s$dGX�KY2hh���&X��~`�m�NV��Ez;`��T����D(B��|��� Wf,V��}Ã���m�8�JĠ��O_c��ʄ�^�8	=g�%���jw�xB���o�J>(���(��O��ϝu��Y���a�w���7M�L����}�c���B�q�E�VM5x��BCq<�5s8L}�
M�_$�t�MW����Ĳ#��s�$�-̴U�����H���?��Qh�lU!Ę�t)x/+;.~�6N��������<��D��CyEAI`L %t��Y���	}>��zh�zPep�{�ab��U��������0���D�����y7K�<��/&s�f�6�"S]뒅9�h-{�sޞ���,a?!��c������M�6��@��˻ �m�x2�N��c寽�n!Y�t)A�d�rUb���29p�'LZ�o�b�$�.�gn�1Sq:����U���vi�Cҫ�WlB��8J��%�o_ $~T�v�VV:ꪈ�E�AU��^����P�C"4���k���R4��7�(�lk+0-�� OT���Bo"�! ��bt��v�����'���^����R�ܨ8�f�V��w�>�_�WоN#�����8�ڗ>�!ak�b��Gjė��1��	�B~�}��mc���҈;�bG�3/��tT�؇�mps8Mu���{�hһ��}���m���~~�	��I����h�tT����MP�d��n��E��!t˟ޚW� �o��^�Dۨ�6sLtH|>��'���]�=�-,�����`�"���^�F.(��HR�<�#�ԉ^�=E�A� !�q�Z��WML�X��I]r�$C���d:�l�c	��g�|[�:�`$�Y4Һ!H��/2155���7b�PfV=r�t�FI��_���0Mú�O�Z��T�*D���S,S�n%f��ߕ�N�!S,Q�fԖaV	1���i�~��,�2}:O�^��<J�J_� ͒��#t`W�g6�t��X���a]��+2O�$yN���5П��$R�#
qLe�R��;��X�|����R3R�qJ���z��ʐ߿O���d:8�/�������������n�>3�U��l���/V�����>�����;]s�dA�d\�;��^MY���?7O�b�������o�B}NLSS,��>-�p�/������_<��
������+V�#�R.��-D�p���E�C q�ŧV�������b=���Äew`艚�M�����8�^\�����J=�>��%	HP|3��`��u��#82n���}�1�f�;ň� _�S��/�p�;�m�NM[�AZ7���Q�S��޷C��f�Jô�!�x.�����U?�v ����+	���\^E;�_���gӎ7<�"{� R�b�u���E���P>VEY3��kb��o*U��)������ԣ��=z�L�F��8��z��8��}K�G__Q�rշ�~.�	�*fegP�w���*�	�G���F�?������ �U���
8�?�i����Ã��2���')᳸�����nK2w��5��MŃ�+��e���Q�����4�j��*�����t~�B��ة��OE��ӥ���a��bG��Ee�I��v2������эG.|��k���q1#��%l�	�z]�^/��x�q�D_�p�'��C���'�t[�=_��OH1T��{�f���6���_ 	�W�t/�+lj�E�b�)�O�M�U��R�'q��b�ը_{��>��dY,P�!�o�I�4�U��{!��N�
��!�o�bt��n�p�D}���zf�Cj�����28`�e�ZW��j�Ӧ"z�ޱɶp!��%��ސ��R[U��RU޵���#�7\�p���_�u������M��a)cp�ɶ�	={���I������;1�T�#:�}CY�3�8���DL6���ѵ���8��۟ZʢЋ�զ����1~Z�\��#�X�ٽ�!��=2�������S|������͓��V�-���o!��Vi�YW�h"&.��A��'8�%r�.Z(�'�����;��I�:F5�gJC�l?��Y�:���~�V8�U)*�d�a�m6���lO(�����:.ݐ��aք*����Q�	v�e����J}�sm�3�\�L(&�D�+��kR���W�Vd��6���P��N�IR��nr-j�e
��6L�W��zU�����x��,ި���f��r:�-n[q�׮Y����|q-�
��Bl�2${]�X�I����+����i�3�9�W�����L�7-��6	�ǡ���A�0/����y���5�����u��ɓhFH��S�I$���S�j����2�"��K|��z!��������	����o~���9-d_#�k��*�?��$J�S�.:<����q��{Ӻ)��E��������J�݋?�-�|K�UpY�����>S�r:��Zd�}%A��	/�g.�O�O3w��(T������e����:�:��w-�4����W�tÇi ��Bc2dJ����K��I-;j<^�.�f�qr���1���|�.�:V+�����+a������B������ �Sñ��~;YSDa��_pÝ:1Eoث1&|��o$�p�%�_l�&Jv�庠�X_��!]O�܎?# G��mԜ��&F���R@Q
ho%�*qCMys��s�$�Š��f�_�l���6spk	�`���Г{�zt�0ѩ�[���,:�W'lAuw���<ҝ�1<_I��(��z�
�)�2�����9B|�,s����ߏ|��6��x�r=5�h�N��;�!��d=1�fuZ��Хj�\G2��:��ܼT����(?b˳�5�KT�J�\.��)j0s�LY�+)�;���z�,O���Y�[")5�f�ˁˉM
���"tGY�˩t�	n����|�Ҷ��*Uh�D\�rwmq��fc��/s���2���x�T1l���Lh��& $d���ȥ0[�'��:~5J"�����������QaB�����Lc�{�QN���S�͝�G��4�cؖܚ��:M��4A���_:0ѯ�������xlq���0��7��K�_�S0��/��G�a�����Q]6�bEd<������s�~ZM���.���}2�j<�拵���LP]��\���7�!rt�tWy;,#9'ᗗ�����)Df��,�@�7J�d����IVwy��׎����~م��ɛ:���%�ŝ����Zoo�޲\���*C,S���-�R+��S�Mx8B���4VlYp�]R	e����6y���	�㛘v���h�$���Q��Yd|Tx_� 4tCv�\����3(S�c���>z��ٰ�+����`��h鱦�#�o��'��ͪ����6b�Yv��7��'��>Nd�Zy�7�w��a�쮃Vp/���.��i��uə~ �u���ۧ?�V����Ǹ�Qhw'�t�ǆ��f�(G�'����h��ʏ�I�=(ēcq�؈��w%ae�0T�J@�]O��V���ڒl~����S���(�Fv�lf>���_F�l���n-l��f"1��|~2Xs�}�B���B�n�xHٿ�H8
�{�rs�j�����o0=�8�{y�����$��k��hUO=b�M����H�C���#�[N0�&�y��+K'������I��Y���5Ob��
�jb�oQ�`A}�-�9������
i�|R,Gg���PK%�:��oLqж���_��a��~$[� �?5��I��GR-	^�oٖ�\Q����{�|�t��jv�ONHt�m]��T�u-��(^�l~�����U0G�5OK/lE��o�KD�$�����
�w�������]�8��
�Ķ����ҝ���&V�$,[@��E�=�Vi|��m9�T�����9�U	�8����s~�G$�d6�Ͱ�[���֬��c��������P�k��v"����j�>�f�$���ĝ7�1�7��y��N4�_��T 6�ϑ�V������q$Rb�?&g�Nr�ˍ�����2�l�aA^�;�C%8�WH�S�,� ���f{�h���ׇ�-�|�@�e�U�5Cjn6����0'cwd�lp&��|,���8����mS!������L��x]�boHi&�mp ^�v�M��/�t�nc��!��4�1bS�u���P�ٲ��"�1z	���Mz�z|De�نv���sb�<y���Zw2���j��-�+hՕ�la%�5����/N:�sL�I�\.�2����ދ�^�������;8��,�y��h�e3����S �WC#�V�`n[nV�_���Q#��> ��1jݥ1�^����q���pD2���	o&�1U����-N����������u0�nɂ���U�0{T�Ki����u6Z;���j�n������<��/$���j�q���W+���}��'��K����x8��ӈ��\ʊ}y5�]<�cȤ1��.D=
�0u!|J3�E�x0�)o8��dؤ6`�h3Y�4\��'Xg�9����Ei��ݺ�:�4����!Snc�n�ܯ��ȋ'�4C±��8���o m7�%�_��$��&�݈�*�ѵg�)����k~��J��^9�<�~͈$�m�+����/�Fؾ�}tYWr��؈���d�Ս�fb�\Cg��Aתp��*W�~'*��d��
�D!^��=���;!Ɋp�ޮ��������7�gv�K;br�>��j���P"�,�.-��*�#fq �N�ĪK�O%+9­��h|��6��r�iߘ2�lZ����$���va�|���8�~a��c�)54[d�s����GJ�̫\�!H(8R٦N��8	�"�v�L�=;�h�D��j~:�دT1�H�#F��~�:d�S�bS��_�����}�^�=q�p�~��y���맼߉�B�����W�Vx��������{XoD�']Ha�����Lk�ԭ!���gj�4����4��P�P������2���f���t�|e�] ������e�P���X���g��Uh#k�@��)���v<@Α#'E)QW�n����<+s�F[h�S!+���lί�û�=��^#_���z�!yS�,A�����?{��Ȉr��lv�;�$�D� L`��ߝ)�As�Ț�Xr��@��T+FW����Y>?�쁆���A�!5b �����'=D���왣s+U��QgE��������$�4&�e-�r������c��Ի\��^��\O��c�o� [��*�yD͝�oe�6�p�N���n5���ʟ���s��q���*#����n�&�ژ�'�p)�=��,ss<�p�<<K�����=��4tak����Cr���������eӲ5G��E$��P��)r��Sņ����ZV�>�[?�ݜ�1�W�2P� ���G����O��w�27�K(�Ǳ��2*jכo<�1W,��9��g�ѩ�c�/��?�2ㇳ���+D��o:�KG�3q#�����ژ���EEl�E"	^KQ��^h�AB!��1���̗�������<�rA�U�G�q���W�6s������:�KL����<���u�io\z3�o�l��i��InM1o��\��alX��MNF��8Qщ��e:����3oDp��#���M(2���e.�L^=���0�b^�Z�H�w�� ����WyɎ�ty���q��uy���l���O>"��{��F˙��S�]��D���\�����R�����m�L(��ct�>< �6CϹ^!%n؅i�X���X�J���wC�,���VV6��x&=z�(�Y�(b�!W�B��"�͙��qmF��0)p�����������yS��.S|�j�5�2M��^Y���ew:b��Mо܌�8��" �\��Н�؃���O5Z��7�oa�ۨ ��S�X�_00�^���3���O��<�74jZ!?�r>^�i�[|U��	'����=}��K/r���-q� qp!��xJ�q�QMi����V?�r��~E�s��m��%�<F}�q�4�!��2�u��4��-�\Y�ndw� �٩)�hn|����7�F�������g4�o�w|6��(�����B���`g�"�@s�J�:�_��A�z��F�	�Q�M4��9�a�O�2�q<@h����X'Ż�|w3����1�Q�!��{7GiP,Il�/n�ٸ��zJ:����LA�!4�C�E��p�H-:1u��h�֝�oL��hMgϺ��;�	-Wu��%��/����V���e����	�կ��<A����t9��#u�kl�'0e.oY8J[�m|oooc�W;��l֭��w�]oX]ﾣ��ff*�l?&<2��^��f)Q *�'�)'�|ct��`3���U-�����ɓ.�9�����5�|VQ�sУ^��w�R����v���9�%q��!É��=�#QQ��uԅ�����}h�^w6\����D�j�U���q}�������D�o=!��cD僻(��@���B���
���xz�0?�~P$�$y:%�y]t�5�9�J��g�����^`顮�o�PZYZ��#Y��Xp�M8�#ލHG���s�c��_4��Cs�q� /��b��ř��Lb"���lAw���SY�5E°���[���P�Ũ�C%i����-/G.̑��MAj>�@����4�{�Ѐ��!�
���]�:W����Y-j͉�))"^���/�yfC�.�PF�O� ��3?�1>���x^���q/5]x��l[�!��[~ѱٟ[LX�D˗w5����-e�cd��1�(
e��\�4ݙ6�#R����u5L�<���L���O]u��9�:��.³^��#;0�(F__?���
�l'����Ob�1�ЕOM6�ǥ��y� ����U����ҁ+�Y��G7��O�)m����sQRHeE��_�^D��z�n���ck�&Z�P��db��Dp�KRf�.�;@��K#��S}���{�w���tT�����!�.=jTƽo�c��+��5�x�7(��/߫���b�\L�>���"�a���A'\]9�k<�RC�|�a�o�X3�ybj�ѷQ9R���;�z&�'�߳����9=��4��Tk7L��P��G�v��o�C��E7N���a���C������ל�қ�g	�!���jZ��gIY\b�/o��<���WO��p��N=F.f�H:,�-y�2+�&}��J0>�'E@v�>!~����I~f�x|�k�E�@�R9�Ӣ%�|g� OX,b#�	P�9������m���̺p�t�R��"-V1�Xy@NE�kNv%��?����=�ͽ"����xv;	St���Z{�Џ��"u�GZ����LeS�YG�֠@wꇪ�d6x��=7�hb�Fgc"�����D$;���l=�G�_��_��;�'�o����v*��TQ��B:T�g����|�����?c�yT�żo���d�.wb3�Y����_r�%�3�X�d���ψC�xQ��?�AE$�3.A����Q˖�J"2~Fڮ�V�
��CJZ�����y��,>�\�>��Ul���*Zl�2I��[N��m�͆�Z,?�����Rhb�����|��g�#{}��eR��{�HA�����d����*�-с>�|#�#艿�E
'
��ɔ�^Y�R��o�?�Z������ ⡄����	}����M����5?���[��*��ąK
@��N�Ekj놎]K9����-��}_>�m����7��ן���mԜd���>f����f�K��q������0��I�oVg��1(B�f���B�|I+���^�_?���6����G�6��}���o��")C�e_Ry ^�~A���޷��N�BK`XN��T$1-į?M�N5,Vd0rC�M��X�To�����p[2@��8v"�ڣٛ�m�C%�s�M��T# $ە�z��j���@��EmM]6��\�h��� �oG!	L��4_m����8��ɳ;�}�я�ő�O's"��}� ���e�'��&@�t�	k%�FĀ	yj�R�8sǢ�׵�gF��8n�;X�̢�o��8:k��bY���-'�4ǝ���[�_�x���tar���*T!EE��k�V9��
��̬�1��qC�K�؈��wae�%9����H	�_��ﰤҥa�a��;���KX?.r�Jj�T�:6n�"$t���5�����w�GP��dha �PfSq�t
��U$�����r�"�4��kq��HG����Y�;�Z`�4�N����
T/�E1Qk�2�#��]8M��C�:1H��]ԟ�*����E�H,��On�f��M|6����]4g��^gɚoQ+���#�<�Q��=�E�׾g�n>���_[�)�
%Ao��Ur�&^�_��_/"4�Sp`�a��huQ�`���`�S)܌��l������w}��
�V��p�|�Q���$"�<�O��]���s�`�ۂ�8��jP�'����k� ���.|)]]_Wc��	�/��.!Vǉ�q�{Xޣe�7�W�Ǯ�K���ž����?>Y|��ph�Y�p`G��B��C�^w���׏x关x��z'�P{yQQ�^F/SR���n!�e\�vʡ��⽂w7-��`&\�G��)��Z[?�Ƭ��<=Y��_��6���>�kJ�X�Ǽ]��t��7;�u��EZ���鞇�y�˞����|�-;�'�f���4�	ޜg��K��v	i�k���^�W4uЊ�)	f�y���="BTwz��?
��N+�q\ڦ���m�!I��A���:��ڝ�T�.^�a�t��XBn��\u���u߫���rv�ߦP�5�_�6Q0X\��7*�_~z��[sy�.�ZiC����-�>� _������%���ӎ����� p�"����-+��p=[������e�}[0//�|U}7`eE��$@��=�a��wR�[������As�{��{7ɔݕ4��yT��<�#�j����������5�u�t�O��J^���C�
f��$F��0�V�M�L�l�O���lӶTS�
��������ǛS��{��qꚻ�6�0�3ڢ��N����F�@:���ZH��ԷG8~�n��A�!3V�M�J�%06rm����ƚ��D��B�v��I�=dPp1s%$�d���ޮG�%wֱ��x>�6�?A��A���[�z]O�T�ǼN�1U]ތK��cR;ߒ�؅��D���\;��_,���r�,���x�٭�hj�)��K���^������n��ү��G��`g��i��z�&6��b�0�9���_(D˴�i띡�{l��5�6�r��kl)+�u9Xؾ��Zj���v֟�8,�R?p˒5l�2v�F����Q�߻�N�˰E��O��DR���ĠU�@�^�G*���d��҉�>6�(g%�!ApP4����xzVQ(�ᗄ�4(8�F<8�3�S��(|Qȼ��"��%�z����V[���B#Yډ }Z����Y�u�^D�ڈHU���P�RA��ǯvK��>�.��@�?�}/�5\m����A�Sgkv1�m���>P�R7�K�� ݄���;:^�Ŗa'vQ%�6^��=��R0�|�V�P&_U��������%�D"Gb����b�%��Y��}�.o���k�U�����Od�ȦAv�)��×�4���2�v|�̵�t�uI��gq�+D�:`�� Q�z)-��j���-�GiP��WNY�
��1�.Y�:n&=̎�]?ߩ��������`�j���V�<_tŞ�65�d�3mx�W8�G%d�
�՗������o�2�b��i���K��Z���m��^�������E�{�6b���E�Ƕ��{�����5�X�u�����i��T�jkkY<�L���d�����a�A v(jѫ>4�����a���;`ei�;_M��V}i��Î/�Q�.���2Q^l�H�Ã�����u���AO<����ݍ`�1�~6H��{���l����3�K�9|��̤M-��q�1�CB.c��������N�S��
A�.}�|�s�(��k&L��J� m	�Lg��]��ep��>��OQ
�=0��٨�d� �No��A
u$%��߸0ՠq�PB��x;*vv�[�F��^�?���4��?�@)�F)�b����G�����'���p (����,`�c�����1�Ր����כ�*���A���nn{ㄺ�A��[=�>K�7���D}�tx8B�csI�;���%s�8d�J� 1	��F��~�x�,�����Е��C��������kA��0'V��ts�.Q��
9�z�eźJkfK���.�hyby�}�m>;��y>�g1T���+ag[�K�'�����Z��g/�����qwoW.��0�-���(8'g��n7Q�v r���=���FK�q�i]BbM�r ��p�\�V���).�k��-�Z҄ZKҦ�/l-j��Ŋ���~��Β��o�`!$���8�j�W#����\�1��A[Ԭ���""* �l�ǩ���in֜�Z����|�F�p�ƋI�u4l{1K��p�(P)���kS��{���f����Rw�dJ`�Ύ껵?�Dq\�
�T;#V�s� �8m~�"�p��@��y�&�+d*�}EI��i�J�v�����sRZ�3ϳ�*����+A�2�tX�<��% 5I�c��]��J\F����q���jd�/)W������I�։J(Zpշ��}o��V��d+F6��ep��K� Q�qς}'��ϾN��	5��,[7����#�q)s5K;;��&\�5=�n�7^_w��
�s�W��b�Ji�%�u�����vLQk{���+_�k?�q�= �&#�4&��+����C����.ˏ�@Y��U��#��z���(��|�6#Bݗ�����Z��rS�JHȬr�~��������6�T�z�&�zi��;ޖQ�d�g�O�[Pn�|x�����'�0����xx�3�auK\��rQUhd���ճÞ0�`]�hС+�d-��L��ǆ���`�F�v�V�I6��N{�+|�֮���U���U����z�2#�)��魊$��d]UygfQ��FYLwZq"�����ׁl�D�K�H��d�-+��ѝ��|�:���5VŇ��PS���y����`_�r�y�k��BT�F�gk�}���ԆF4�(NM8Gi��}X����Ub�9��H�?9B�n�������rb�/p�d�� t�ϲ���,��GJ�#Ӌ4�m+&nL.ˤ�*R�ë��_ya�_p7r���n8)|E|�p�,��5���(��z�)���uXvL}{����/�����[����暛r�*�5_���_�"���n�KS�;��K�}o0����Q�����vO�1e����n蕋�+���8�hK)�	������uU�	uh�`jތ�m�R�r�a+1������Wb�>�ٚ$��Wj�3�PFGZQ��.���d�2yy��M�c����d�DZ��{ˠ8��[4��www�w� ��!�w�����@plpww���έs�Nչ?�jj����ٽ{�^=5��:�\�3w޷�ܓu��!���<�[�x ��]g�@��=W�A��3h���đE3bY��`���_���ßŅ�ʕ��=��puO_��H���K�G�=IB|g%�L�A{>[[ ��'{��^���v���)�~�b���:y�]�b�'�BGh�f����~�ȫ�Af� �=�����a�����>j��)�{���sk�1y1�dh��G�Y^%
q���2�<-J�[�,���7�Y���
�D���+C���)����� }�"2믄Ml����Iis=�Q��݃�6P�]��2��!��S�@���u���qa\w�0K�B� j��P�C���[=B���6��R����fˁ��ܤ�_Uc��C�!�tJ�}T�a���T3B�����@�~�*l���@��ȃ��?� �rl�Efa�;��@h�06���oD���I�~���h�y����xZb�o��br=���wP�8aNA��
���ƧkY���
B��t�JV�����Va�+:ɘ<��
��5�x���~�C�h�z�X	A��n�cT:�C�8�<�b��l�mj�~[7Y`?܆JɤG�:�"�4Z镻����N_`e�K)�k�j:�p��,�.���~���(�71�3C�K���oa��}���K��Z�J�W�)ṝ��1׾��)2�ChSLE���'�������F��K3j�7`�C��/f�"
�~�������������c�nL�Hʴ��~�><���J-w�I*F^䰹��k�2�Ij(Y�K8���X��s�U����$�W��6�!-������=-?ɘA�Q��8)�����_�����$%��qv?��p�S�~�F���xl��0�~T�jY4��D���rx�X���E�	����	�-�/�	�����9(�R!@��V-�y��NgkMÜK��Y��Q
���k���	(��\:KVj?���}�,V���,UZ[�(����!ZY2�s��O���i�~�&х|1�y+���
t���suI�s��ެ>�F��.@�+���{�S2!�7�� d�;/ւ�*� vy��g1B�}5 Չ2�e`ט6���K-����6g��
Yt��9��Vh��b��Dyݿ<���2�/���Jz;Ylpl�C�;�����}B0m��)�[��Q[�ܶ1�k&����Φ�f`�pBȴ�I�Y��c�(;��J�6��g&��Xo�Z!��$A�c�d��x�h�my��6��W�[���,�>e��t?���_~���J��Cp�%���[�����2R6:��y�S��\u�o����������~4���*v���UM���G�V�v8�����k�u�oc'w��_u�_��xH����Uڼ���4�#�v{3���U�r��V��T�r�ž���B�	�T�nA�]�|w���d���M��+z�XP6µ�JP�7�Y����]p��Bx���-'w0�6�=��w/pcP��Bf;u���gZL�u�-�[[[,�0N`�_�Łd[ΰ��$�0W3}q2:��!zXS�}m��<�Ň�d
��!��qi�q�NPdd;��p�=$#�96\��y�����C4L#"bbѣ�0��:\J�$�I+Z<��� aoM����s�Nm2}����׸�܅�C�� :���E���0a�'��,=�H�-���� J�A��?}�D_�-�RR$�O�q��2���t�:�;�Nb|i#�hVw�lݧ�^3�xYjH��x���ᯮ����Ö'������Ó+����-~I2���m��'�a�*�ha�
=<��O2*)���1H���6�ځʖ[��)D��Vva+��π8�3ǿIv��D����w�c�f,�~⢻�N���v�P�ys�b�=��(��nd�	��/����y�'�b<͋:0�`�P�W2&;�s_j�C��v3H�z;��j3���B�����&$�r����p�t#�V�\���,���U�ɤ�Z��@T1ߘԣ��_��r�#U �� |4�y@��ޢ�v���Z��w���0�{�d��v��x1Fx|�ӷ.�d"}���'�4v#T/"��L�9j<�ҁ@L��3�P��ѹ�ڊ΂<V�|;2<�0��]Ќ3�U�6U_��⫱����1|8@YS&ZBS���K��	���bhce 6��W[�������%�?=�e;W�\9J��x����h�G𑸞,�B�1ݬ�q�����96�����֙-~��IG�r8�����|����s�؛y�ޘ���k�JT�q���3	�t�2����g1�OD尠왦Ƨ���fƂ�=�����*vB��k�a�n�S�=g��N8ב|='0���vW]x�xY��ãP'�4U�g��8i�³���qA��tH��{�8�D��u�Ʉ�^2�q�����D����1�4�r�Ւ���J���mեΔe8N�S`�=����M�"�<��E��S���B������Nw����G)�AB�*߇�'/4�ᠼHd�N7}m��d�R��t�W�St�8tn�A�A�n��<�d�5D�8�޿&���6���ORe���͓�c�jzJ���F.-�;��|��k�_�Wi�i8E�������S�3��sR�I��:�Z�P�oQn���Zw��#d�;����e����7},�2��\����e��G���Ŝ���;d`ϝ���Tӿ!/Z�z������汛�I�VE�s��'VYc?ԧ��B��M�ڸ�|X��8{�)�����<P�Ѧ r<���p|\�?v��u��/>�rL�\�g&�?r�bį�/�ۄoU�������y�ⷞe��ӗ��^����"��7�-p������-vP���=�K�\e�g�|;��K�D*�I�C]�K)cߦ8jR!��v����fĸʔ������*kv	��K�N�p��*� %�ל1/�rC�4��y�t�oc;�5 �u[R��M�ZQ��R-~�}�_3���<�^�>Y_1Ru�[�����f��Үh���}��h@��'�o�>���:���ŁC�8�)�>1��38 [���wph-S���;~@�C2ʥ����Ć�V�$�% 
J���"^��o�ϣX6<��!��R[�L�_�`��{Ha��.�g#e��㙬�y���_������ ����Ň@g+ct����x��Op��+D��+�imm-?>�R�6N�pw�G6y�e�e�:�s2��D�r� +	No�2u
�>TPru}on�`J�ĸ�-J�6�H�)Rf�F�'�����ޱU���q��9T�s�h*�H�!�����P8F���o����:cԇV%�8ح��X�]�c�v�:���h2�K9rݜ�+V�U�2j2�k�� �4 �������y9���ȴc����p�,vu\������!�}��Z��G�-���`�*�{<�ݐ�|��!U�����R�Ks�Г�n��䈹(��nw�'�����>�E73J4��������b/O	�-�Ǽ�i���A����]x��D�E	-�[��j�G4�z��U��P=1�����(ci�y"��V;EB�v7!T��&Z Ճt��aa1,q�}O^���~�����͚:��J54�.S��s&g-�.ܑ^�f��sk�d�!Ϙā�~�Cu��qr+�3�Ӵ�I@w��1n�1��aj���ۡ���.��X����]�M�d��������Y[�P�87[���X�z��t�p����{M��YH)�� K���R�-Y�q��ծ�'eZT���)��@��� 3(���ib�'{z��}(���*c ��`�;d����;s�~MW��G�F�������
���`q�+C:g��[���Q��ﷅ7ї�~]F4��[���#�����T1�zi�:��O���=.{Y䈸�C.�8W�TBp�qC���MMܒ�����X�`Q��*tT������d����� U��N��#��;5�)�Ӷ���?5�[5>�+RS{p���LK��_,�z�d0��9����T��u�˝��a��?���ml�)��*�6���uyJ3��!�Qwq��afW�����Y? 4Qw4�2�&^�G�#k�c�ʟYd�����9C�h:Hu�I�uc���bq�u��襬DO4H��rE�'�d�l����#�,Օ�V�l�9CjU~��ulů3�d5ND��0(�2�-����V�l�w<𸸳�B17]Hr�:4[4�W�ǈ"��rx�{ /ö��:ڬ$�a���?6)�0;��gY��x�����A�o�$�gd���{���Qnq{C���Z�on�Ƴ-^�;D�FE�^GG+���E}L�C&�y��=�`�E��$���#��G�xr~����QG�ۋ���AC�����dy���}�X���+���<���%�����
Sǯz��f��'�7@!d��7D\��ܚ����Ħ["���|��5[JA^R��-��2���]:/�Ҏ~!� �2��p���I����D=uc.?��pR�W�y�1���|�O�*M��|�u�v	f`%dG���\t���	B��,������|di�5jzM�~|��cí�I���n����
H�s[������g�xwk�W�ki��~���+83&�����e��
������[(?�_-Q�(�p|˓����$^�<��Q��~}{���͗�xd�Ȕ�΁=�z��'�����\{r�i0�Ra� 0�����q�p؅!��~�L��n�Ϳ�1aWw�852yzz����A�S.L,���O��,�hy�`�t^����!���m��®Y�W���Wfx<1Q�#�xOh��I��+��p��鶌�Z���n��/j��('k�����У_=kSK���[��nO6�1�TD3X����B\��c����.P%]5�.+ёt+ѴTW+%5(���K������x�i�d�ZWt4vKP@��q���׆�e�wg��Ch���)�|
�������5g�5s�wS�c~i��Պ%2`gd���LD��`����Z��LM�����}v�.C�\����]���iIr7��s�'���j������^��b�j�ٯ�w��ٙi��sU�H��d�p><8�TǴ����|S�EE�xx{��h��J��w���y��g�M��}�'��p�����<�#G�<G����v�o�>Y.z*S�bJ�S���-�7�W�UcDP�(.8��L������"����R����fMR#]��JQ�p�!�]�։忪���.��x@��}�-��1�o��Ʈ���%ZK��Nj�+ᩛ	���8��@�*f�����as�p�%����Z���U��o*#l��������FH�q2�֩i����?6��Iqfj;�M��^��к����DJ��F�͛rs���*S�ۦ����h�4���_H��L/�����Ӣ�_��	;-�E|� cw�̤��������%C���Ɵ�w��M��R��J.����oK.�[�X��FS�P�z|%=I������Y���\�_;���L�%!�q_�����8Х�U��`�����l8f\N:r` L�V�o|���V�>B�S�X�UF٘���#A�l�嘞���:��ȋ>/\|��̙_a�JQ��SW
��D��)�Yr���m P��@���P��|��T�y��t)QCsB
��<?�CC p���A���-�W9��r2���+Y�=�SAXl:���R�����ab|�(�x�2�HVǓ��[�b�;F�r��NV��Ί��`�8�8��_���i�`|1\�I��F��K�׌�ٸe�EnK�����m�a@�v3������W�c<�Q�l��vH�R�@yx�AWwn�{EV�\�y�(:�?#HAK1��|3�+6*���Í��b� �Ǩ������&n��u����b�`��;�w97�|m���4O8�~���f��9m��\��?�*����[��m�\���[�T��m��x!���g�&13,��Cg�v�����⸌�KAZs�0���9 (Ef�[b��]��Ӎ�ș�5Z�]��|	ݰ|	�2j���ny��9�/p�ἦ��0Z�)Mt�d�+x����s�W[M� �B���%Zk�s
��CpZh��)o�,�KE��:�ki)�[��n"�0�U���UT��3��m�hşH����3$��q�]�:��.��4��ڷ&y����q{�-E�)�(��S
ډǢ:�-��需_�b����!T�2�,�D��&������G��\h��(lI����	~讥'��E��YVM�ݠ�	񬁭Fő���f�4��ԍN��/�>#xfE�FP�~���d��e��3�z����Q��wK�
�6����L�.��ቹ�ng~1�e�"�өARm�z�À&Lg���:�؊j����/�
��3�Y�I#k'NߩF���f�L�=��i��L.��z���?��tyq�d�6��ʌa�A���>���Q�/�j���T�Z<RB3î��N7-��������ݠ��H�ۤJ)Ա�'�95���u���shʶ����ՠs�*'`~P��<W�1m�QDf2�D�Q=��V�-�Z��g��G2�tR��./b=�~jr�ɫ�2��I��k'F�Sg�[�Id�to��|	��iB[�a&St���S$>7)
+�*o��Xs�`�|wqϚ�����^�q��å+�p\�5i�����$�ܢ���:\t=l�\�|73��b���6Ę6���ԙ|�s���m��j�#$�U.ر����>Mp���e�G}e�n�7����m����;�8nC��a>�3jZ����<����@�ݶ7���t�#$ R��fmq G�㎲�M�����uZ˖��������!m��@�^���։�O����4H/bվ����
���li'��;�;�є�����`�R�%��Q���e/���pppk ���aK~~�6��E���A�_����Nˆ�@�j��թ�9���E�3����ڥ�¢�����^d�I�9оY,���U�h�drݩ�/�e�9{�.����	�#[a��Ŭ�N���U��HDd��L�t�rY	m��d�S	��FGER��Y���l�jEz|n�'<�͗�5����WJ�ͺTO8������/���Jǅ��S�0��œ��r�|RӰ�:��c}�zfj��HA���曇�2�C��J'n-RbjYu4MR�UD˓_,��ki�Q�>9z�֌�-k�qA[anlP �Ti�	�@�*�T���n�2��t�0x���'#�s���`��DI��3�����}���o� t���v�	�P����g3#�XiB �6>�ݹ��/���sV�9�XAI��h�CX:ܰ�����:[�8�Rw��,�������Oh~��y{jÇ��t�ĸ�vd�a�w1D��t~�p:B���2\T"�K3��E}7�6���t0��mq���}S
�/i w�uy+#�&����������dF[)��./�������h���9���o���s�&1�	�JT�Ќ�%��K`�� ގ���&��?�l�H$J�tC���u�vy�#�*?~�u�E��5�'���;�b:^_�w�����a���7b4}���_9�����>H�{z�BDl2Gp�@��M���3xf;;�܇�����&�-�2����u �6��DL�
`�3H��^�,�/�W�LЈBkn��L����鯲x��l�\:�~m}�	��e�H��D'C�`�Ί�xM�3�-a{%E=r�D�	]��:pK���	���j��Kj4A��G�/�S�?��L��X���rA�5�LҔ��I��5w���&�E�B)�� �+lO��m�"�]ۇ�9Z��Ձ�ܒ��>�9�2����7�aJ�-ƽW��j�˞���qp3���>y��.[���c�\i}f�wd�'���Y��^䔙��qkb�L�@5�#>X��'����['N�,T��8���oI�'�H��߸j��	�֛�)/���ys`ܗ?R~k�X�
�z6��X�~Z)t�jza@��8��D��Ù�e
Ң�9qR�Dii��\�wo�n���b@؟ 6�ʙ�)���@�!����~���f=�"������ #"t�E����E����|�(���
�L��3Ol2�@����\�ɟ��"^��
^�@9�_�����o,�d�o�K�"�/���d�ԑ���KN]�d�؄�H��X�'-�z|	$���S1��~��&%%�P� :���Z^�+fp���7?	� 	����\����uL+.!Q�L��,��h��Eq�hoeE�a+�?�m��'sny7?CA�pE�םSS�):�"	R�/)����܌�[B�ڎ���bg%^�(�X#e�;E<�2ީR�]�~��Z�}���T
�(�O�V�Y)y�P�
_�m���f[i6L�;%�g����Z@ҙTH|!���%�
7�!� �o��
|H V���ԏml�a��%��;M�����$�cDt�=�3��<o^Ð������sVa�!��+@�޽Z:�9=J-%����;#��>8B�ר�|�gٖ���1�&"��`{'���z��MJU(,�п����4Z2��W�����7w'��~�7���{��� �)�nW����#�}{y X�tWZG��1�F�(HK�����w��g��}毱�ܸ̰�)��d�u)b�Z�Ԯ:݉�\/\}J�9e�ꈹ<eQ������5(�_��a�ǆ���4������d�FV���PLVG����TI��� T�����כ)��`��?X�]|4�f띞�5�� ���w��u���S������:��D�>��,���N����<�����GFy9���	 �s��r�c5r�ƿa�8�µ��=Y<4��HL�"܀y���r,\_d$U�_��Q$�A�?����xq�43G|Zf��Q��{zQ���R���W���Y��t����b��q���@m��ݩ����Q	����@�3�d肂���*���	DN��v��p�6ԛ�H(� �V�O�6(����>��A�R���A�c��-�L����u�j�]��E��_�8�S.��f��������5k����*)X�D��Z;����x�(F�Ҩ�J���mkm-���{�p���Osb%�e��s�hd3!���$�u�
������p�kms��V<�ySNdb!��	�x,��cT�3�����aߞŐ�Z�eTPL��8P}����E�2�N��N�Y���9#&�ř�1�������s)���T�@c]Dk�Vh��R|( @�5>�b�T2�n�l���U &�f�iV&Z��*�>d�v���ad��G�W:4Y��f���j6�|�Be�<����ϊx8~W����?wD!i�R؀'H��=m�n)ɊrYi��%�6*��v<��W0k���r^�<����4�v�	�?yq�+�r*V��K0����0�M�˺���n����j�g?�=C��F�������5Y���V�n#���?ǋ�{�
e�۩�>r8/c˭J}w��n�"U��|کg� �&��*�dK(<5�����o��סT�ѹ���h�/^;�u]����Q�X*���2�V�v�l�A��������D������.��X�ڱ��4���x=���:F�Vf�-9�],�y���$�ʬڦ~XoAVk92��(�%B6�h���o�]'�nD�!:&=v\��0�j;�`�]���*e�����,<������Ҭ���zAݔ�qR���T>��:�nfa)�<��\�i�:l��� �9B���|O��ö�T�$�V��� ���T9��G|��f�nH���Q�Sl'�8W��#�r�pL}���%q�(s2;������o�
�:\��x\"��]�9;O�NKqN�F�VP4��()VX�V6�T-�X����ْ�S�Q=���G�^������u@Ӧ���f9yQ�����AZ�ޓA��2����Fe�4P�o���Va����		��]�FD�ʲ5�ro�W}X!�;�i$|�ؘ&ֶ�ܥy�4��'��S�v�+3#�郎��W�����~2���8��FW�acl�V2z��h�w�E�`�+|'��M�����/�a�܈��^7������I�'���a;1��wn	d^7��~W��ie�ѣu�V�s,[x�\�x#�?��.�m��*��WE()��>Y<
.T_�gb�F��q�\�0��J�ό۲���|�rS�(>5b�R^1�SW���5F�ps ��i�3��30T/�pa��dPlμ7�?���M���?�-����:��=<_�����$]Uɋ��:�v�}	�3 фW'�l��.�����sJ��YO��Wm��'^;e�-�9��r\�ܶ�}�W����[W������#��HL���5`��DŲЇ�\�O�2�PO��Z�E���9�"T���\`���}�����tE$tŏ@�!?Y
u��4Bb�
[���<G�4�]=|�>MSF^<LW�z���?�=����
��&
�!��W�O�*N��-{|P`&i���"���Lפj��9x)�b�n��U&�Ĺ�	��#���|Ć0���k�\D�4�*/Qlb�
��-]��S����;	YD8|�F��a�����tS7Ҍ � a����4�u{��v5mE�#�}x Qb�6�N�og�
'f��^�P�wml�6��.`<|ܤR5ɷ[��ʹ��R#�.���@6Rz<���Ǣ�c�����cNk�7��U������y�֎�S��h��p��--��H��A�=G-m�uk�K�X9n]�5�m��ʪ>�~��D>^�3�J޷ �˫��~e��~�}�b.���Ζ�1_I��)��B���c�.��K�	{�L�싘�U�������"<�#|n9VbL����M�ejo���x,x�s��n,�FH`�L��u��B���A���.����
%:��%'H��@���M���d�ٗ=��tj�*{�y`1�	>�t:<P<�l�JЎ�"}���{�8^�xt�a����M��7�
3C:�U���*�D=�Ƭ��*���Գ��(��B��q�����%�VRr���*k�R3 �oth���H������֭�����C�q�9�l���)�;���C�9B��Ȑh5�SG�{8���tњ� �CK+ewS����;b�E�\���A�Gb��Gb��zǭc����\��t[�/Mx�H_WǠ����ޮ7x}��a'�w���zWU'AtS Nhf����l[��ד�l-�U��#����������Jm��0[x>�!UJ�Tx�=�t!�]��HֆP	r���z/��S�,�b]�:D+�Y{��4r9
��֊��	�[3����k��|t��~x��ڟ�<�-_�ۍK��5u�V�8�^;��H�Ŗ��u��
�^�t���>�	3oىd��^(be��54�Ps���tE�@�y��m���T��9)��k�+E��7�\��
�B�:�L�����t�	���+��{M��q�Fw�����B�"�K*	���~ӻg�n{|�Q���Eq�^{ϟ������u]QQ&��������K\���Q=dsws;���L��:U��(0ob*�U�����,\^��z�Y���lt�0qL�?4���+/�-�7����^�4~-�XK~#����F�--����^��H��qga'c{)��D!�$�?�kc]J�])2���S�,Ҝ�aaP�_�n�Y�5�Yߗ�r�ϝ/�|�'h�������˹X ����9���O,F�F	i׉�_ϧw��	����
U�$��F�� �\[l���~vtT�^�3��I�r%mk��R
ʼ�:^i�.%�!�f��!�b;w�Njq@˧˶UT�+�D@=��Ͻ���=��_�!6if��}��hʚs�źKJ�#�j6��B��|&/[|<A㝳�`�oG3����#<N��pm*@�쁄'���
x���:$��Z���8����!�4���{�)c����^!"�;8�Ɲ
������}(��;�_��Ws_,�1����6!O�Muzq��u�J�ip'1�pG(��K@kS�! �؊�=�X����i��EJL���{�De��;-��҅��uY��Y����)a%q=փ�1�J�.���j��w�K��N�]��|�|���y��m	�M�n>��N}����B��U���E����|L
.O�Y%W��,����k����[�(��������QdKq��U^\�M}���)�:�z��	^]ʩ!���Mb-3pE�˴�^A��b��>���v7�w/@�qu�с#��o�6�;{��N�K0�Vb��}c�Q��u��W���f���VdLu�b?M���v������1���^K�-aǍ]��f���Y�y�1݉e���i�L�U���>qd	K���eu�{0?���a�s��M�,C<@y���V�o���Y���f��"N*P2d��$&P�֊�h��q�A�j��KlԿF���"�=��g(�ˏ=;��ߍ�&�<!$bKi"����'.�������h�튍X�<�ԜHi��4� =	L���)����SH°2}���=��ʴ2�6����G�5ѰZ�����M�S�uCxt92O[��\�)7yB�bz����k
��h&�o�lL���4C	0g�d�X���/;m��Z[%���Y����*�T�ƅ{�'�R��.���&��u��R���s��a��h��s0��s?fx� �>�{Ԏ8db����C�Z�(��z"�=[��8��B���*��֪�WOʬN��s��B�3�	���J�8�8����4ژ�˘�R	ܗE�U��(SHԌ���gd�crt��`$�C{�m��T=�tѰ�Q���"�Z,d6�E�Cý�f(e�U�2T$M@�v�w�����M�n�1X�����U����NǠ�vf�<�G�Z�n$>b����ԡ��l�DSa�pCC�P�3cw:���Rc����e�Ϙ<����f-�)�܁?�SmM�ڰ����_�CDYjLS�II��~�Ha��aӉ�@�Y��\�J�tS�i�9����0L���8��y��@-���w�E�1�h��TOX�IS��z3�@�qO����vˠF\;���x�m2F�1����U�qC���k��d�#q��}�`$�=H���<׳�^�䠪�uY�BQA��P��� :�`�S�u*4�.�������x댒�����zߝ_�\VT��}�p������y"���	��������>�`����D5����o���������:Þ��4�ѷ�H	:��a��z�GQRK}k`ݝ��-']���s�)��^�x1nH��w��ùۂa67���+��ŷ6�#jj;��p��o��7��	Φ����t�%̓���nj�ӳP�Z-��@��]y�9N�?}��J�M5�(��	aTH�A�"6#��!�xẌ́�F��$�PYs@�v���w���*R�e����.��W�����Os~@�)E����,�~_�1�L<>��8�,�������J��X���ꪅ���&�Շ���>e���Ea�:bj�È���E������?�N ;���<�t4EP��s����FN=�&x �U(;��.�^Z�D�ѯ���[Z�	B!�*w�Z���7��mMg�%��6%@�yl{�-������S~�^���"�2����3�ٸO�O���N{��27�*���,~ �@F��K����pٔ~��/���B�EK���K�ꙛ�Jt�Ej;�]{
D��bG=��?�"
g��G��Ҭ��}O�P����J�i�����#�����Xr�)vB��s��X6�oI����7j�n�d�O5���f��N��B'�}>^	~�h1j�)7jc���u�މ8ӏ2Y��R�  
b�a�:�.�%V��!�y��xB�E��a��� a��mBllh�X`G�]�㳕I����*[�;,�0z�T�`�dV�:�œ�9�S�|�����}0d>������|��G/jƼ��7ߕ���.�t�nm���O�]��C�Oh�ȡE%/ ������������ͧ�޹ϫ�(��dt��)%9w%�#qu�ؾ���F�??t�����}���/��Lt�
�u�"3m�Pϑ�%��T����q?��[h9�hGS!����2�xl�:r�^c�TUf���}����6��3�	��̫l�=�-b��q�]-n�&X�t� �)�������j�Յ�0�y�sZ�Y0ՏW�糅@S{�ĒW�ko����	�nx\��&�Td^��W���Ρ�g�.6�ˏ�D�H�s����`{��P\ ?k_t�g��J/��J~��˝�m������0�r���X�@�Y�1�j�֜ϺG!��ְo�u�(��3R=C>{>�`�o�|���Z���Uz2%�����^�X�� ���'���+Z=Z`�����tq�0���B���/8BX��qq|��O�~���Bm/�0���Fr�n�3�N�t��"��}�/FRG�AKD����s�3�|@�fzHh�7�W[�]r��w�������}u��}?��֬hЙ������&ȧ3����j5~�Mᵋ0�R� ]��˝��c����(kjR�:C랆�ӡ�9�@k9JRy�o�?�M�6/,u8Z�R�v�����ܞZ>wE@:��H'��S���b*a�'s��:�;Ĵy>pi�$���d�e��Z*�S�:e.�ȷ� �/�0f>(SN�EV8��a��;L���$7��+����P�3�Ƿ;|A�^\���(�<�e�=	�1U�;�G�!�V��]/a�%��N=��/КR�R��}ρ�@3��,�O?����oUm�'�:vkv�[���J��-��^'���%�x_���w�Ƨ)D��#l��r���N�yr��8>\oKc��$~H^սdđ6�����b���3H��ƽ>�:TIC�&:��{5��O��Q8��$���`��������%%$oA~�d<�B,�t�ܶ���=�?�<iK)xC��A��9�S���z�J��j�2��O���G1p�}]�-öʜ�e��j�ֺf[�Z^/��_���
d�(�4�r�PJ7tu9#K������*jmկ�'e�i~�*W�ɠ؉-;�r,:,�,l��$N�Ծ~�^��e?��F�'�`��i*�6����r�'�,���Lif������s���2u(u����1�i Mm�S�θQ墣 m���~f�]�g�뿃 �(ֆ�7�ڕ\~!�g)F��I�T?Z����S�xJ&2jB�h8�Z㬽�d�i���O���D��yS�$�:�]�X��'w���!�e���#��˴�*�'`��7A��53����k[���F��ڰ
��������h���ˢۜ'opv l�B=�c���8z�E����K�Sf/�_b�&��J���߯I��
 ���>7{cs�gIK�h�^Ղ0XFA�Չ�A�q�3/p7y��<j�^p��U%���R�2��RH��K��1&����>��m�	��-*����D�w�y����OZF�I�'�/�|RI��n��33!��f`�c�s�`A{D6�U��p2��Ji��+:s_�oc+����6�� @���h�xIY|ˡ_�41�Ě���8t��׳k�o�,����,4���W�4Vp})���b����P���.Qnr��	CI�r�v{�� ��ބ��f�Q�uB�s�T�[��]�/s0.��D���)����p3��=F�$n���_��K��y7(�]��B��>5���u��gx�Zu_~���H���O�Ɓ�,w��cl;��f�����.��qg�j��(�c���6� ��[ ̧Cc��t���)�%Ά����t�[��[����5�Vah��ݣ�b��޿��_)�����w����xg��9�b�8��R'}z������� y��={�� �M�}�W`&V�B�d3 U�_���$j�����4�~�v���'<'�T-��A��xd҆=$rY���Ch;��4�m˖϶wi ���Ѫ���Bܵ�b�� ��>X��P�Hk�"�1���q�ʍL���X�ϭ�|d
�*@\��[�k��h����VR�4^
�����y_�"����X]J&����8�f�q+w�]��l��%E���e/�%7�����n���͎0��8;&��K����G��թ@���[u������ ���)'*���&��f�fVun=�Њ
�����܏����;�k�]�|��y����3�
�W�$��������+h�Lpw	n�.Np�݂������sqww����0���5��Z�0�������ڻjױ��{ֹ�t�������x���B��ƫ�����}�_�%n�Ų����ۀ����Ҍ���G`Buk�43ݹ&��+�ڷ��ڽB���Α��}�bY���8�$�9_n��$xܭW��i.�����m��,���qH���U����d!.#�ï��]�s�9���Z���5S�H'�!#U��l]wZ����]�$V:IQ�M���z�n)�dG��ȀS�6��Y`j>e8�&�;�Ѿ>^��|(�Z�ݎ,���R��N��i�{�;ᕈ�V�U�l� e�N�i&Ad��\�u����C�?�㰃��k�Vm�Ϋ�9�
����O�~�E����~PYE��F#� {�1����u�����������l�Y�.����i>�Z
��yg����(���4�f|\�3کk]�lJzVH	�z�s���<o��{c�c���;$�a�u�j\Ҩ*U�L���k�md`=��j{�¶���	c`	�A�������{ډz��s9o��Ͱ�yc04EU:��S�*��A�A�z�����~!غ�)����1�䮇fB�"�x�ѽ�}�'1>�-�����v��8=1���Gco�gF��AZ>�EH����='+���q��"���\{}&�c;�",�w�L9����QXe�6v���2E?��b-���_t�$��"s�?�vÞ̹:,ȅR6��C{t����9q����l_��f7ȉ�7U4���=��fۘ����\��»Q0�1�8��Ю���0�J ��������%^ýkʯ� �r�Iu��uW��Ic���wk�s�h[	�4	g�w�^�������8���.��8)��?g�(�<�_@�~�����M3�����)^�z8����AP��s����
��	����Z�pl,���|Bp�2��wWn��+z�݅ug-�A���5Ԭ��%�[�sB_�6��R�8T���jA��OuH�eƀl�8���FD6�	����z1������R/�^����;s�{y�K��4H�c�9����F�6͛q�!�IQ�^�(ڙ+��C��0�����M{�K\@��,uԶ#�. ,0�`���C�4g�y%K��H�=wC��0�Ú����*w׬!ܟ�����AnJg����I}S�����i�o|I_�{gu��QC�0\�����Np�ϛV`Χj��E�ҏ�a�|y3S��u��Y��"s�e'=�;n}&����9�2��[�8NW�ڤ���0SO��݆O��.=|�D���6 5���c%&Ժ'=}إ�U���ҕ�O���V�����C���t/K�:�W�S�N�hVF�!�K�QĥŮ������̾�_3r7��wٝ�q�����u�3S����i�u�)F�)����>�-D���B�,ME���S�sZg4G׃Sv���l��l�x��P������t f�;~ ��bH�6��J*V����0�e�4�f^`�ڠ���}+�y���f���n?�xp�u���1��χ��ǖ�@�kT�َx��ni��%���>1r����s�c��<b>��m�61�Kܠbq+�n�����O�VF���Җ_�Xh,U�2����r[G�Rk:||���.�-gՂ;S�`�ǆ��k��;.a���k�a�t\<�#����ם�*W̻��%V��" /Sk���i�snU�԰ż����2����ёҷ��*����,F-&l�� e xwy�01TD؇�_m�K������،~q-Ҭz�l�p���a����5�Y?T��(�s�Z� ����{��y�&��.�g$XI'1p;ּ�JE��IB��D���Z�|�u���(t�w/G��J*����vGD�^��T��0���p����ji�k�,�09?��5�g��;�)�.=���*��� ]`S�S��]%)~J;��}^�~�(�S	%���G�摤c��Jmw�t��t����G,{>����K�5��;��!R��_�ȶi;+4� �+�Z�NB qg��ּJ�ui+ |ek,GQ�ޝw�����h��n�0g�v�T.w���rs�>
�V'�۹�E�l�� '��Q�
V,N���U��`�EԽe<����L����Ի�!t�Ƽ/Ѳz�0)w���}�CAL�V9F_W1Z+
F)�*��0n���}��yht�&�y��ƪH�������N�#��*փ�C]l��pT���*�hǔ��/?J?��u�������6��E��8��~}���3r;�nu=8���iA���ob��ԑc����q,����C�L�Q��<�"�N���������H����gւ@,��L'Ʋ� �<���)V	M�R�%�/�)A�2�a��ȝ�Pݙ�����y�S�؉>>	]?X����\�l.��=�u�>�0Mw�p���-����dr
�BE_M����s�]�o�Y�[-;�ܥt����ܳ�Э�U���H9�qiY�ڄ]R^V�f۝�%�7!��	0a��%_m�5j<Q�4��+:R{��,]�S}.�U�n�O��Q@?\�@+��F&���6|.�Ƴ����?̝���Z�&�Tյ�#�pO�.�9��e��rQR{�A��'y}פKq16��
DB%D��t��d�XJ�I�ul���J����)�ص�� m������v«��D���<���R��r�/�鶀���*�3v�V����H0��6�՗���ޓ��Y�����oA���f�f���6^��G����kj�}�~�O���!�G�8$r���$�x�^v���^�T�7�XY�E��4Օ�����)�PtAگ�2.�n���y�W�K�%�uy���v{�(�̇R''#*1��[+<��Niu���%K&ZP9~�=�;��s��4B�!�.C��R���.'��-)HSBz�u�e�I���A����g((�K}�Lų�g����E��V��osՁ)͂��!�i��%G�W3\����n��Kع�u�6��k��蛡H.Q�Q�>��\�l���� 8�/�K�/�L�,�)f��,sB��YyZ����@(��R�x�R}}��LM������HH�
���UnΫN�ap�ӿPb�tK�O�&_?��S0�n*��8�?X�FR=��ٳ��ھ��!ޠ���}�&/Y��T�y���������=�?(3/�G�=/.4w�? ����/��6�~ù?|��V���p��[m[��Ȣ��j��EqX�c7��Y	6�W���J<J�SZ�Q�(��1��!��r�k�c�w���S�䞉 '��;�Z��3D[�Kъj�n�JS�����#�3k
Bs�|t�)�r��s]=��S��1��$��#�d7������i��3V��n��pj2BWmP�s� 5$T�nXV����;�r�������iE����o*g�	���1�2��&���x�?B#z蒭)�^`e/�5d1�*�FGsJr�w�]�m�'�����&��8A9ˀ��]ES����Y5�tU���=:	�c��(�ؿ�F�ڪ�"��i�����J��d�H斔v����Tg�Zc��[��� Ϥ�VIFrz������"�]���R�ѥ"D��>��H���E�9 ��d����k7ڕ���t�^����'����PB�@������ؔ�;`g�,�8�ƓC\���|t��UQf�E�ː�f��֘{Y*q�*t�<����M���ѭrJ��i�R6��Ps䃉��r�t����w,\����oӰU��a�����oA�)�{�%�?�>P;>{,�O��3,�6���,/br�f�GNd�Ќ�+�$����RGp�D*�;�Q��O�1�E�j���a�Ʀk��'6ս��w)�������=a����êW|�n�;B~�`�,B"|ҭ�K��m�)V��O�p��
��r4~}M͐�7�Y@���E��zjQ/^����;T����9�oo?N�U���&ew`�HG���1A.Q��I��cc�
J�t�ɪ lP-�YvE=�J��k賐�"ҵL�^�,WMUHQJ�����}��!��q
7t�����0����V�����o�?��:<�f�"�+���#}b���H1г�� ��W7�f}��$CcW���>N����< �p��}(��9���ɚ�S�K�/'�!���8�rVV�ྒྷ#�+#d��O��<�-����K&����j�wm�ۆ|��F�=�>�]�����C��O�'}}}5��4���b0D`��۵�:$(Z�6c� �j�p�L���������3�����������2��q��3j�X�Q�����&jkC�����Y�� ���C
i��U;��v��1���֤�H�<n٘�T�����a��1($$?7���J�6''g�+:��p9D��H����ϟ����w8L������YeA��:.�I"Z�&Ώ���`n՞�������a���-�Й0p�V{
�K|S�=�k�CC���5!�fN�bn�S�GC��pxoow����7������&H_�?��e������Ē����ԛ����o~<�.Vi���ة��C:��,�|NKK�ҥ�������}Ɵ�"\"� �֌����2�[�<�ި�րC����2V�����$��j9O#�Ń��C�]\������E�Ύm�q�O^X�ӊ�t45X�ZQ�qg��v;�~X�9H�g�ebd��z� j��)T�% �u9��E�^m�����=���������
W �q�{�E����� �ѱ0������-P��뮋(=h��y��tk�s�����3{TX��rI>0��z���(�8�eL)�	8Q�ׯ�{�_NJV��b�WW�Ηk!-,,R���t=�w��t�L�?���l4X$����^4�t���˶y�:��Sn�uѩ+ңT_e��6�����K��P|�J�QgK�����$qt�N��3��8�ڔj��Z���4[�ɼ�	쬭���FEC~����8 �����Qы.�twvv�q5��'��~Q��)���.�\��i7�	ä6��K�h�z�of:ǹN�����?[��&�An�6@ϲ��p��K{X|�{�$FHDV���6`�3Ĩ9h�H�l��`n�*,��̾�<��@+Ms�;�e0����\��Z����i�3g��?���� ���(���*wo,ZM8��c\��P����Po3n�r��A�3ێu�xa�7}���{�ީ�B���ۆ�S�Э�aX�W�پ�
�a���p{�s�>��^i�	�Bں��~O�?��&%w2�g��N۸q��̂��vx-�ج���L_��o3���~��Mu�����c�V��&@+��Zct�i�3<�{{rX�8�z����TSv���\�9���i ���{���^�ކ��Q�#��j�[�8���yj����~q��&�#�qV��W���F��L�s쵘cGj[����?��'�߼Ħe/ʌG-��d�O������|ן2����Ki-���桼�-��a�^���G���553�7��Q�yB��H�����L�l֚X⨶�X|^�P�1n�����H7�/K�eU�[5��(Uc���xs���wB}yM<�em���Et�}�AAy���-�`=�쎻)��Ά,�-NL�{�zӨ�/՝�wZ�����g�!��c"@���gv[�e�m�="F������B<T���eI�z���̐�n��Pe�31T{`~~F��p���y�t��
����`��
*Pawӂ[�{�J�ɻ9vj2�SΜ\-y48�[�zF�ӱ{��_����Xv�/�v�E�����,JmX�&w���e���xBv��受�+�~����,$'����нJ��B��A����l�����erώ���T�e�3_L� eߙ��._h4�'=��MP�4)$���]��S~2����֍7O�k����J�xIX��P�D]����������>�!���yF^�����@����Ǜ����';VB� /�@��Piv�GN��>�ݮ8䘛_7&?O0�cO�H�o�א�N��:I5�%{�sVEy�����H`���ZxS@�R��R[���p�֨aT���&��5Ƶ��@�:M���5�9�Jj�]IBn��:OC��h��71@��-8��)u�Z��G,S�M�Z��W���G]��[��x���S����[�]�O����Z��l�3��5��7띖Z*@�Z��Z_p���As+:h�쯗�yTX�?m�=�4E�,�����ѿJR �\����*�UM��I6g~ږ5��A�/��^Mm���2VA�R�!��q�z��}�kzF>��G2V�[��5�t��=���~�E��I:;V� �%+-ߺ��u����cp�s��۽\�c4��$��9wф��O���F�gY�oxz�7�[DZI�B\�P �.�;�}�
�����*�k�nwvX�1�,G��ɤy˙n�w���Ȉ�V�	�>�� ҽ�}��w��J�"TU���:�8\B8�j�rX�?�\|��p��w;""��X�T9�5>`j3�m.=���C�˻����VT�XH�+)O�.iG?]v�K����Yi6 �n�EfW��~�lC!�ɢ_+�S��R�lq |����[Cԯ�=�u{n�gN��s^�7�d��f�Z!a����R�^��^�������������Zҵ������k*�ŌIAGx^���P`'���p�+?Tv~uU7pWWf���:S�Bغ������tX�2�=���t��&<�������,��|[��4��%ԙ8�k�����׸;��p��-�uݝT#�﬍DIJU "@9xs�cRf� ��B��9Џ���(�ꆿ
a�w�VV{��i�1��i�<�ibg��f�go}F9���1*2������x�c����r5	�y�y�x3e���3'�t��X��v��~h�@<�����!�|W�IZ)s��@i�KOޚD��������f?�*Tp�z����<�8�=��\k<��.,��L�Ǆ��p����R3�;ι¼�'�!>./��,[���u�a���tȚߺ�oS��s��M��8Pc���g ���|���ZYCfS����(��"E5e�mCȈ�}%��E�}��� JU(�䔱�&��P���d�� �*e�h����Gu�u�t�+kl�E�L�y��!���9!���`�/e�̡��y�U��X��l��_�M�4�v?QmDt���2c�Ldsӧ	�W�j����"��b F�#4�_|n'%R�Z��	�M�Oh`٣���\��=2��t�"���n:o���iF��1�����$/�=���;��@\n)pu7�PT�$�y� �������^>(1�ĔCP{��z��HI�u��{�G�Ę�����]��������1�X;���MU)�ZZ�B)���%YJk�Gb�N��	y�����<��]�(E-ɒ�R^� ����x��)N_\�J�Ɓ^�ݴbi�Y��k��n2���l6�[�R�_x|_C�=�ŉ3k�eKSYE=�m��G� �������E�ƚ٣��?�'d
L0����m"���Æ�/�E�9)�:B�z�����b���P���9���^������)P�	� �G��r8�[Я9уy��U��6c��QM��� Ր��p˻.G��{-�x�>-6TG��O���Fo�đܺX��[<[�S��$�#��z�ܚ5=�\Ҁt����&Zd=آm��rK���G*��}�c���\��:�Wf�p�/}��p˼ص|��>�@��ts6��Ix	o0��i�Z���'��^���z~ �͡������0{��s:i����~w_�-�a8���@�yJr�}�H���{�H�a)�Hw:#J��/�K��Q�b�~8��_�.�5�i�c&*H7wn��?��%�kS������ל�2��e:Q�.q��� ��U{��p�[��߳�}��G��?��~U�(��+p�̲�<r���IK����4R���\�[
�I��)n�p�Ѹ�S<��Ԍ���W���8���0�iz�@�����%X�
�xޣ���-jЙA7�ɼC������h��D����tЭ+�6�Ϭ*42�ݒX�F�~��>gˎO����P&�]w{�`�.?��,���Kk�b�_^:VZq����z�&�«=:,6��?�X�7ɂ�(�3y�Ģ�gl]���pFۈ�<��1'��N�?{x!t��Ҩ�Ъ�V��:��2�MWq���-��gs�<a$%��"�����(�6��*���=��,��1>6����XsB�ޖ7>��N*�������M�z`�p���Ǒ<Gm�OA��Va�&6ӻ<�'�~{.³���f�[����el�&t.�I��F��5��<�r�,�n�c�|K��>X�/�����/�	ł����kh Xn���]Cг��C*L���Pl���a5���T!� 7j#ǟ��J���ϾX�g�%��<J���*c��o�����B��[U�!~ޭ�-�,���P��!P������`~�^�w���/��	Y�q�Y)�ҚR�����9�Zz[9�T�#��_��I��3N���@ʧisE�F�ñ� ����5o��X���8c�\�\`����~�D���Sx�����חxn7��ڧ��t�֜l��SG�_��ԛ�j{\^:�����9�{�t}l�[/j*���~h;�I�0�{o�6r9A��뀭�g��5u�=�Pt�gШ�ڙ|���R�OV�~\	oV�]7t;a[FK�qz��
�	>%�5EE7���3O�;r�>Z�X�N�Z,��V��߄�Em��S�R6���*���N����f�f��u��n��� a��m�ʋr{���-�ݯ�7�A�EA�����������!-��Y݃�a��[V\�B��&����mE������:�&t����u~,���A3�" ��j��Or��{�3�-�JB��w�u�<&��:b��ýo�߉*\s�ER}�پlq	�7�B�[͔xau}�&�}�y�y2����~�a%ê#��a���y5�����&6K�"�S��a��fW�J_D�ϡ�ӗ�`�e���0��uø���L0��l����g7Y�R<�hAwy�[�{����7�	Wm{\���m��[;��k�^��$���"�u���Q)�<Ϝ�����P�aO������y���T9�YB��o�'�	e�l~OW�.�G����5Y_��`���P�u���շ7o=�ʰ؃����?D�/{E�T�WҜ�9�Z�锫���z�'#t^y����r���� �Vg*��Ap58F֓�]��Q׻i���P5�;SmhJҾ�\�<��g	�Ӧid�7����dK�\��Pr�ԗ	_4����髋��ݽ�?��9�ʱ&�o�󗝊G�+�%Ǜ&�[]��w�Ni��7E����F��A~�ْK���P x4���}���x��W2c�.���3���������˛^�U
��BF&�,b���2�|�rf.���/�)�@�UiX��nʔ�.��?������7��Z���GKk׋�iֺf&[}�����;��?gX���D�N�[:X6� I�xF�������eK����ۀP/#5;JqW��D�5
�����E��}� [1.��ߪ�G���_Gؙ�t����b&g��n~84K�m�89.��5/2�1͇��L��3�G��G�jqV�\��]�tvcA��0��^h�F��qF;�}������a2(��$�%�������%o��|�p�R�O��țoFq��|�f�({���E���Ƒ��a��*n�L���;�yہ ��]��R(��3.����s��"�2����YB@�8j"�?%�y��h��l��t?�Y��>b�N���7�s ~�Ei@��`��R��U��V�)��j4���x�R,�#[6f��)E!k�(�0���.��W����kF�Z��1���9������>�IZ���^߰ )�&���Aݙ]�--�2`��>kM�BMf��$.���N�>��a?�8�	c���~Q|��h�8PS��0N�#~�f����Dm.j����h�+�7����i��[�ܭB`�F�|P�c�7�x��Ln�Ӂy��@��
Y��_�N��k���%~� �My��j��%�j �^?aO�������~���|����iZ.��白���V� ���Z���{2n���Q�{|�xMz��~E��'�c�̀D�ѯ��ޛ�r�A�k��74v������h.=a�g�`��������7��~�{�`��I����(��E�>�+b`�%��4�do��������޶漱�am9����ꇸ�d���ms��Ru���m���[��8�r_d|%\��!��%�HY�)��5ӈ�������@�:��']�O%�����N���u�yi~%�؉>Ƞ��5�u�yj��p�bI���U�8ש%����������'G�8��N�2�[���y}t�K������q�w�OE�>.�h�F��*��i�)O�L���n9I����xi�i��F~먵�R��^7d-��u������jtf�3.�!��&���M���⅙Y�s������W-W�ӨX���(������O1*��l��1�V��`��fG�fNcNO��#я��}�{������K��4y��r�����~�6�i������0�v���f��\|�� -gQ�2;b:��,�JY�V����
a�In�mȒ:*EJ:YD5β�|�\T*��d�V�-��o��x����ǲP�ܡs�U�9V��h<��xЯ6^D:aP�p��U�����0�{�X����+���7pu�*c�6���2���٬m�u����	��LyM��Φ��&d$���փi��R��o�g��j%�,S��P寶y���պ��]�
53]&�N��: iLx�ڔ�Ζ�o�;�$G��F��e�ǰc�Û�V��S�0Τ;��Z�a&Anj�KYV��|X����i;�_w����>�b\�+Vki�ב�K�=�q��>>v�mȬߐ�Q�MM���f�s�ID�^�~�H�/�l7ڷ[�k@=�Ǭ�?���ɪWܿ�U�����K����"��k��N��b5H"��/W��v�}�[�9K,� �INA�y�d���k���ʊFL��#�тg�G�O�Pbm��Z�\][�_!�_���fZ��P�=R���Nm���/�D����(ɡT���.�_����ŗ�y�v�jI/
?���1ٕ�p����n���z,}���3�&�-��f^8���l�#������(� ���G��S��kZA0�z��"��}�$�:ܹ�'*��R��=��E=6�5H�˝`�����u K*�1n��U��#rI����s��sO�3�?Y2[��=�K�#6ĴNQ�<���#��1:r��k@Ç�Z��N�Q�����w��Ύ�a�[�E�nҳ"����u����?�]����,�i�偑:+-GNG�AF�ߍ�/�� ��ѷ�xTf qn��m wb�e�MC�}X�R ��,3/'rQgqm��")\�CPiyfw����e>:�bo���.�m�q�0�i4P��Q�D˱���(�}��0
��S�Ǚ��>VV�ƪ{T�'v̶�m/��_3��>�IEIG�����x��4Z���(�@�4�59�Y��)��r#��n퇜��M�����8m�|;">�B�tI�*h�'��N$9��#3=2�
Uv=�s�y����0Qf<�1��p!V2}�#�F��8�p!���Ud��r��^�vG�8����H������V��r�Yeb�� rw��Qs�1���F�����%����5��k.��o��|��b��K5�ꏒ��ӟ�g�V�Ȝ�{ŦL>��_<����7��7�F��H?��'�z�F�ok���PFvy�)�����,%�ۮX� ���y3ЛH,�ܘi���6��n}P�[�L�2b�����L��B����*n��?�?=X�\��n*q^q���e'o'�PԷ ��@7*�Y C`e�8Y,M�b1y�Tg�|bS�H�oŋig�B<^8Y�Q�^�J���j�g�����ݜ�j�R�Y��Q�a�K�f;+�z�y���jg�����,G�U��W������@��N��Zz�/��Z�TK�(&�k��-���cO��^�e�>S^�o��A�ɹh�f��<07�}?��r������䇚�0	9K�Mv�!���%�Z�`e�����EDE�-��x��$��$���)�7W�nD����#���&�Db�nz�}/z���\��\����ƍ��r��erd�=�kˈb-�Ž����^����3%���AE�f`����6	��Љ����A�mRY��I� ���e=J%Q����~�wv�P�5\� �Ap��tJ;���I!{trI@��Ek��Qu��;��_�Mv���v��T$��͊�B@q0��l�@���5٠��Nro�ͷq�z��q�غ��X�>��QK��Wf�i�JDb���1�K?�U �<[SϹi[׈�fǋvrR����/?��������#5j�fr�r�בD)Q���,d��`���'�����+a���?��ӟ�{�:	�VP.:z-W�g'��U
M�$G64����vٹ�bMj���B�u���%Ύ��vH�vP*��ԁI��rP�iл�p<J����b�,C#�s�"�م�9r��Q��B*|�:�h�a�կ�j�1U��iqV¸��[0��4�/��*@/�'�+���C���~�J���Q}�v��b��W&i�F�ݰ{� �l9#���@V]S[+r�"RcuGhl��#��\���ʯ�&Cv:3�� ����k?��0=>_o(5�����@�CV�E6��a�l7��S�������?!G��i��J�]J�����դ8.�/���-$_�g!���i#!r@���N�$�FM�Kr����������fZ���[߱7�G	�V�5��F�Iޔ�N!}�)'�n��ǝk� ��V�0��*D�Ux=X6�:m\���[�CGl��vo�}vb1�|�E�.Gϩ���+e�{E.1�a�
����|*�y\h�����FQ���T����Q!�9#�?VS }c��F�z ��NԆ���|t�����7P����87Q�W����i�zO�I4���|�n1D9�y�e��|�,��;$%����cn�:N�@Ԩ���q:ǧ>�Ν�ͩj|��:BT_+��
��57�i�,g:>�f�Cv�x�{F��k=_�y(G�O���� ��ҥ``�Lc��g���aF��C�;v��N�<�Yl�b��\]���Z�;�֑�R�j��=U�C	[e�U�ٗr�߿���	�Sw~(�r�Ng��)W|�$zf��]R��S;�s$������F���w�Lm5�P�rp�]��g��(�R���,��$'���|D�!y�g�	��(����j�Ϗ�(���Mv�!���#�\���m�P���q��-��'޻Ӛ=�N+����V��@Y�M���;��ʴY}[�XrS)t����Z�5���ݫp�l�<��Iկ�<�&G�㼼����
�fK��	$�-�
|��o������2�xFط4C�J_��&{�����M�N�T���V'/�J�`���k�B��	F�ҸEslSѯV,-�c@�D��Pl��|V5��Q7�94h��#K�	Zo��Fw�g�G�� \�<�Exp��mI����0#��A�<����	7����i22���owՙ_�7+��_^#W�L�(M���u�c��r=���5D�"���ٝ@�F@��������|���k�A��'�[Z�'�I�Nr�P�{.4D�j �K�2�C�����'��(�T�\%&��J�g9]�~��jv;u��8сv��F��V[MW�;�f�R�M1T3�6R���r9��8[���=�#�4���!��O:�A9Cd��W�1��A~��Ģ�>nϑE��瀍�K~�P�
���ު����=!���/�Y�?6B����efaWC���]`�wK>�E���ռ*9�]�\(��|��Ւ%,��S�}H���Iw��-���%O7+�K�[A�2��vAT���sS�AqL]e���KΣ &�nm�K��)*D9����	3��v୓���:�������zO=C�e{̿��/#�6��h���)ُ�=�9�n��Њ?F)~�,�I)�=*|��f�v�����M��BE=J��4�����̵I���6A�����R�0���uH�4�~V�z�c�6
�_U"[~D��~
���O�-�2�:���&i.kS�|�B�
�0J&(��@)KxD�T/-6|*$��,~�+��MC����³'��Z�[���Š/�Ք -�F�5�r���g�Y�����J�,��-ݶB�G��DV ������֨�4�Yf��I-����Jl�F�a%�WQA�R��3�S�:�[�.ob�N����eSހ˜��=v��3��V��˳��lY� S��4 �0������x:�r~&vF�/[�������t#֍�
��j�]x��9O*#�
Uπ\o&W��������2�<�3Æ�9����i˶�
�	����j�v�dn��K�F�W���:�V��D��e��#G����X����;sy�n�#��E{~�T-����K��FmdIi�Ə�Qш���>+��8���6��UL�AiHV�q(�2�j�<���J1��ó.�D��׃q�t��k����7�<�l�&��n�̎"9l�Vq\�lRHWZ�}�M�"t�/�$����C��V!�r>LG]i�	�Tǰ��=rF�r���l�={�u1��g����3N�'��,��#��N��%����u�E�(�%��*���-�ôL+�[x=�������np��.�6������=�U��r����z���id/�8��s�lY� ��8k/^�%�#6����f3��$��LdL�k M�06K��s�]
�1�|[.KQ�9����s�IG8��7�s��$���$�AX�9�K�Y���@�=#����ν� ����m'������<�w�f�3�>d���a��E��>��U
zc{�o��̱����v��%n9X�٧piGG~��G(�:���L���п0��ċ�3�hX��(ҳGh��D5xj�'��<�C%��V]���A�������둰!<|�n� '�
���"��&���W5����!�i��_�Bт�M��� �hw�o�J������.�E˂
�HQ�'��ȫ^_���Ul��F�?>5"ok�.�E=n_B?-YU�E2U��iwE�ph_�Ȇ�M%4�Tg	���1�0M>@�Z�D}v�F�O���#�J�v6��E�'t?�
|Z6W�[ME�5�(�va%�÷��%��{�:"�#��o7b�V����#$���[�����A:��Z�ɉ�cT�� 
c���aG���K4RJf�8L�e����r���+eI�eʽ ���N���A�����f�����m��t۩t�γ�R��!���L%\yD�V ��*������/xN4��NØ�R��nm��@��2��!m��>R���EC��`R�㻩!��+�����j��k�_o?���-���4�J,�t�o�l�`��H�p�/	j��CD�y��ίԔ���l�ߘZ]�P�}S��F ������J���ܴ�`RP��v�J\����|-��?Q
�A�él�>��6��T�[�z|�-������j�k�>I��/K�o��IA@7�|��p�m�r9P��f㆟�:M㞺p�PU�l��*���e<�����V���D���Ff��.'�MM�}�����i�q�<���4��,>Cz1����YE�\�_U:���'U�q9"f�G	�1r`H�V~7-�N��2�g�"��;k�/����V��uX}�Lk��Rw��Mr�obЋ<���jZA�s<���_E�g�2�=d��8���D�Rs;���/)�0���%����A2�v0�N��� N|�%rs]\���Fs�v��A�.&o�N��ŦR.����qΕ��T�V��u�(�ш�Rl�Y�f\�v�Sq!M�3v8l̈<ig���Tg!�_�$���������
�-]�L(�GP���F��KC���I&-��ɭ�@O�m]�,�P޾!��=I�T�޺��v�����
 ����[��̮u����H��{ڟ�`�PǇ�˝��Ҳ�\y�:����*��v�z����������l�ֹ�zW�wƘ�I
��p;8���I�OP�Ty��XB|4�nǳ��^#t!�t�	O�LW��1�¾��L�Fz���V�ÆHPl��@D9J�.M�aκ�/�GZfÑXN_C�`p�l�gn���	������yU���Ǒ	�X~�	#'�EabOl�3�۾���k�j��e}�hH��阗Op��i�>�*�R��B�2��vdU1��	yPO���4�M��O���W�(�Xh!v+�D��M�B�l�^w��+��Ο���-c��K��T�d�i�7Ҁiu謂B����3�5LFq7e��xr��.�1��Re|��YnnEX�8�zjj2�%�!>�%�^��p�!Ŋ$�Xa�%'���Ȼ C���9{.��+�!�6�ۺD�ˇVh�w��j���ޟ���.����x0���N7z���o��(��k�������w	xp�";�!$ƖE�o��7�Z��e�J��U�wC۰�2��6���Y����.Y-jU`���K��WQ�3<�l1$"ׄ���P�ߢ�����;Ap6_sĵ;����]k
�(��;�>r$��������YC�bM)���B�)k����`�4*�f^/S�U�J+Ą��Չuޒ��E�x�����2�ք���m0�jy���O*J�O���$0���Xޛ�Q�إ��k�9�:�Vp����
G���d�H�������D�i�)��Rn�t�Y($�7�����8��a�4�Y^jg@��_K����J9��[GvS��]J�g��[&�Zq��~;��Y���o������h���-�B�t������x�z_k+����?�/Ii���#}����F@�]�N~�Ss,}���Z��E�p,.��!M�^.���p�Ő��gdf"�]�� E�4<���?ԝ��9�.���vh�?������99K�8�b�H;>1'��k�,ʗ
z    IEND�B`�PK   ��X(	��I�  &�  /   images/9311ee57-74f3-4b31-a8d5-48402682b362.png|�uP[�6�'8Žhq'8�R�����=@��ŋS�xq��bŝ ���M���~�����̙̜9g/����<k���"��M�  p�߼�  �P䵂���#����Â��w �^���Oe^ � �W/�<3�31Ԟ�]ݷ�=8��36�X�g���r6��de��O�ɡ'z�����ל���f1�.��
���E��q�\�ѡV����?�m�_���\��g6J"J �o��x�z(��+��	�p�����������訯at��:�����<3*�����0���B��U>~?9�%�# ]["2�c;�^���5��6��n�Ba�|��A���1(h�]�I����qaAbO4����^��7=Bcuv�&ۑY(�zL�$���\úҋފ����2/i�K,�>�����-���р;�����(m^�@@ c�?������8����`9F/W� g�~��se0���A�
���m��� (m�8)���||�o0]M1�_UZ�{dD�����p�;��cy�O��&2Ouc�k}�r��A�F~�s-p
B�� �oO���j߈F2�1�b���>q�i<A��N��ZC��7;�FE��⇕h����š�#� .�6����s���x=(�r{ǽ�-�P��
k��������>��k��e�ܔR�%F����+*
��0�Ȟ<W�琍��E,nsc�r'0]���^p��d��mvL-W��+'D5�W����3�"�H����O9�H�$:�qw2�-Sl��b�B[����E�LNO�����h�WÅ}Ӟ�vL��=:v|�k��������II$����_Hk�O�+�Gh{�_e�������i:>e��\�+4J��+��,�f�Gr,Xa�.���z;;u�/��4<:t�[���T�����n#5�aUN�ι0����B� WW��qqq�l��
T�󘬆�&:��X�꼁���9b���T6�Wts8}F�/v�A��X��У˃7�s��87w�.��L��Y! �`��f�PO,�/����L	�s�˦�Z3ӌ�w�=�F^�Z�yX�g<��ɱ���!�+9F1z�"�I�8���M�� \���
5��C��,��ÆÓ��w���<�_?����S���~S1
-�ΈH�Bw��R������7��,�s[Z��:�0K@i�bb��u�CG�1���(B8C�#���|��BE���:��X���ڔF����r��� ���'	�"���.W݋	գ����g�����$�'qs-��#%�p��^��h��C,��(���!�][�z���J�[3	��6���vʑ�\�)��=����w����8���'��m�C������B������D�8L�@B����!o�n��!E� �nq���4���7lzzz����%�����o�����Q�e.|5݃$�}�r;� j�&[k�}���Z�Lw|:��iV�����;��������+23A\Ibc���~�9����~��40�l~5K|/y��e��X�K5}}���ɤ���{���b�45���|)���+�T�N*�JTO��R`L�������o}0NC�:-"5��n�rDd�|O7�s��أW�����u��z����u?�Ʉ�׃�C�Fv��&	��|���{:q/tS�����]�E-�j_hA�[#�G����Z��T�}.9Ͻ]\�Z<=�H�W��K�aE}��W`�-g�Ӌ7�P��`�P��fI��?�6Wkf6�e~7�
�/s��LW�{��J��kX�)����K�x�ֲ��$W&99yr/�&(��lhh�9������&g�c�+5�_SQ�@�Ҏ�u�NVu���-oPEj]�tL�=]^�T�Qu:lg�/�`~{շq Q1�B+��@�,�GFb.n
�Ӌg�JI��CW�AP���
T�ꥊ lI%�"��9���q���2Md�Q9�Ln��h�N��)_M s�U�q��z�z��җ�f;	)zU��I�<��>����ˮ�PPTH<�9�6�S�Q�a1٬R�����E�4
�1���y����~A����[� ��$b����|q�3QTBP�p-�g�	[�_ff�9:��^X���P�{c�`�$� S�˗��GA��=���&��y��csTc��2I��Vz��xUs�wg�(�h�ԗ�3r�K,�ON�o|���ߎyE�� �-�[��/�6qU���Ui���zag�/��x�u��:�)���7���O�4��H�� ��_o���*�f�gJ�	��'�v��ZOd�_pPP���З<!�����)���RŢ�bΘ�~��L��J�7������~�����9`�~�4�c��sx;��eǘ!��d	t�xC(v}����e7���7&$O�����{����H,���BA@E�\�e_LA�����m����P�'�v��Q����w��VL�`�A�U����=�t�H�Q��5t���MV�� h)�#��An�Q��h��YB��7kIh��V����[+��ދ�-���Je��~�T��TR5
��ձ�mYRb�����%?�y'����,LC%�(��F��ы!��m����C�+
�(<�w/�4^!���5�O�yI�����u.�v�yG�Ԣ�/K�]����/�4S��٨4���v�^��V�C�w��###���?��m�FJ��5��w�'f<j. Ӎw培��WU�*��8)h^]�L�StC d��7e���7%^�E^	�v[V�[x���;�+,�������l{å����s �%8:75=�͍���L�i�ozϏ~lbɯ�/� Dni��\��I�C�hġ4��L'�A�эZ��@�b�J%���/.�b콺}FJ�50H���5�1����-+�^oE�t	?��T��Ce@f��0��?M�֤z�,gGm�[�i��Z?w��4��B�d�Wj	[�v�u��y����@N���d���js���J�j���	�[����6�rc���T[����$ಓc1�w�h:b����*:�w�dg��0�ԏ]�<�^{�_|�3g6��#^6<J���b7(�F��Y��&6ev�-<����7
�Mו���)�[7ېa�Ҧ@��o�,��_F����ռcx^R�6u�'0M�%$�5�搕 0�Ć��Ļ.6��f��o�\RH�BZ|�����`���=&t�(}~���K��K6d�b!��8�<Rxf'XхJ�|��9��h�v��W���t5����T����}�����}	(��Ii��wR��(p�/�V����"{3���M��+;2D*p��TT;ו�M^ޠU�F�Cf�Zr3߈�Ӳ*&��}�_�+G(ۧ�0�߂�Hc\ r4(���uG㗝L(N�w>���F�D:��؋��ӛ�z�IN���̜�/]�W�&�'�!�~�� �W�o���c]�;8�Db	o?H�Tp}��'��8��{���"OI!4����_���'����Mg9��-�ѝ����Av�sxhwV�1�5'�5^���v�R�����\�ZW�J��_xdw���H������s.CaaT�C"�+��9H���p�����dT�p�J����q�X;��5��'��c�����mw�h�C�jKK��1�����ld���~��x~~��b��w;Tķ����V�Ë��[.�!%k�q�B��~�Qm�~�#gD��ѽ�`�`>,-�΢��r�@�6�����{�v����'��7��o)��GDt~�����ݬ/�&.!A&)ݸœ��|���g��W�w�)ł~g���P-�C"�h�_�P,��S`E)Ӕ������}L�����)z�ž�H��(����|*X�
��}О���N�w���FgҚq4����ɷ�P;Ko//uR�f�*A�P��W�5֣�J�J�3aϟH��t���,�c��b@'W�{�\��ٝ��IO���[�٪ђb:�����Z����A&���ք��N?�m��7y ��'=R�g|�*z:��e�d���B���Jt�\�5���|��V�$�^���p�n��p>[\;w���b�`�C�2&����s V�������!�%3okJ
�RF�M�����lU�~��. �Ϣq#u^��rONj��_�U?j\F�:9����+�6�.��Q�2�ѓU�����g�ѲZ�t,�|�{CfK(F�Q�Sе~�����,?�-�(�'|ΗT,`7;+m�̦��O����j��8)**�s�k�5C'��z���A�,�ZXZ6��
ܬ��9>�>ggϏ��z�@�0���1+�`�ZW|s���\���[5�8�XjqDhT�4� ϑ
b�W9��H�F�F���i�8
 ��VWӄ6tϛ�� e�b�� �-�T�ʦ��Ю��*T�pn�rqN��.R�)|O�B�0pg���CX`,}�m�������b���'�9�C�#��M z��_�N]��>�8���AK�b6o�	��KY4:,�\��҅����e7H�1h�xm�'��/�$�^ �ߜ^�w)۹��8`y�0��A�-g"\��7�P����r��OZ��b�P�b��̂
$�I���b
���9�d(y���QQ�������A��,��B"�C�q����fig�&�J�1b&bĻ�S���m.�{��Y�?�sZH+��}�����VPP@R�՗�(��	
 ��譴�{�]�o�Ч�(�W�;�cѯiO�j͂Q!�5���������;j&&�~�?U
KY}V$�����m��-�k<h�v�Y�5b��tP�����L\v�s�7� ����N���_�NNN�@O�1�T^s �	7h�뛫���/���뷰�]:ɔ �u�RK�'T@>=�S�6,R3�D��K+r��h9&5�1<���FFeB��[�1͝��-���g��i� ��f̡s&С�<��.�%K ����pm�#ݷ�7cYu�}�R��c;
���;��t|�~hw`��?	��LH��{#�S|#BpK+���䠟���}�Ԁ�G�&��<�ha��'1mz������c��PSa���=Ay�Q��=�<���N�R���i1�XR�شݠ��ӋTK�G�h�f��D'5�����vҏT���[I�\�gfcD\���e��*�8_�٬�G��ue�cr��:��C�t�*�Ă7��^��< �z��߿�UUU}=%��c��mk0b��vL��/��#�W[��S7��&�3/��T�&G�
�c��m��:R��Cb�M���2<_5��c mݹ��tQm4~|UP�̮�C1ք�lSh�6�Z�1�Z�6�瘻x0I��A�5��������s���T�m_D%�]z��?f��h�U#�꒒�����F�n�:)�i��� �Y�	�d��q��9-C�V�5Ԃ�����..tZ	4r�����c�#���'��!W�� �
C���2��2��<�50�"N�羹LUR�t��N1C�+Or��>��+��@�O�nF�/N9��ȩC�h`ˑ���ʎ��9��糎W��� !<X^[�6�С8��M�[�q.[j��	���7�!�
'�6��C�Ǳ�֩ۼh��q݊X����D���Dz�����#�(=�0*|�z�u|�VUj�о㥧u�%������SP`�{�D�B2��01qW3 ��5SV:Z��W��yы]��r���50[��A�A����ُFL�Iv��s���r���t$�A�2@���53C)A���lI
l<R�������ִ�;!J�ݲm�B��fe{�q'�`~���Y���︬����T���0�?!�o�8���������b�|�wq�Ɋ���~����c�;�'�o���dO�"(�pӎP�>�_���g�+�̈́���g��ZIm}?sDU�|�Hk5�brk���S/���<W��;������.%��ET1��l>E�I�v��DA��3���1y��x����T@��^�mt^z���0:�Vb��h��(�;P��]b��Vy��,�)伷�I�1�6y��IR�c�m`�� nSq��Ħ"ә�Z�;����"�&�9���7#X!�*�i���FOJ2(+�a��kp���Ȝl���)�H2d����$y3��xR���F�N��h�������k���p��̓�2?H�/�f��=�WS�̖A^�/~�6Z�6�Y�]W ��m��K��	F5�����Z��b�����X�Dm��'��Z=�;?>2Lp�ay͒Z �uɤ�m���f����i��Sȣ��Q� v��vf#�%{tI�����YQڰ���D(B��������o�^�Gw�Sh)���	��ި�O���Z�M����k�N�����@�`��;�cB05��SO�=�6��5�*5Y���(���8'ъ��@���l3����KL�E\��W��<�'Mdr��*x`d��@;b�NS||S~����U֦��x�m��u�%a������қC��R�-Q;�͡�pqJ2��L����Emj���sy���D���l�����zK�6�Z�]c�����Zy�ئv��i�,e��Q����ɠ�!�q�α_R:����^��v��{���W�ul���^~~I��&ϓ���>0\KAA2S� eu\{NIt����&L�����5,X�)_^N�����;�.����������5c�ލ]s�"��ȋ���-V꿚H�u?��j�?=p�����Ǝ�v�~���
ә�sdC �����w��\��=��`ѱ^��yG�]$MN ��7[P�v��_�n�NƂ.ā(S�<�Yn��@쉊v��MV��1>A�s
���8PvzY��W��b��t�^|2���|.�I�
e�]A�!�t��^�Q�N��]C���6�*h�6\k�z[;K��sPE��C������@1�?�ڨ��ī�x�.�HMl/k�����kQjĶ��H'e�I�@����q������]�;�X �ݒV��x��Oq?|�#��U��!�%�0�
i�����}�����Xx�����P��LX��S�\��cL�GEX#��w:��������t�_�������~���R��aZ�|�w RW��j�3�#��S�3zU�94_�k�ӛ�d����?⼢䑨�Ju��P��8O�l$�.G1�Ky=\R����t�
��dB�RA(���"4�Q�J��1�Kl]A������+��֯ʰۂ���y�Obb�9V8����K�V�_�S�.Z�r�w8�"
�VH���+r�n����9Qn/	sN�[�H�����Դ!-����5=���AL2!�� �t~J����ͨo��2n:���^lTd��9����j�N�Ę���.N��6ć�����x�Fl����H0}m�l)d˭B-2����j>i����八�0�{ukԾ 0�+���{����Ov��r2�.d��A}]�n�"s�n5%�l4�ǚV�+�6F@}�=�
Ȯ����=����R�g"b�5<2π�_����� ]5L�ژ�HȈ_�E|[˂	V#?� �]���|�f	m��Сu7�!���h�[)Z/OL�rn�� �4
�f�;���)���zg�C�ww� ���@P�<���t����,��eK�1���~)����5H��tMI��a������8g�=$ @&:o�o�6���1�/�`T�,�B��0�l��[x�
j�yz,���)2�5s߰����4g�:`#H�}7��Xf�?#��oRv���'�]���U`" ;�G�hic�O%�_�wq�M��]���T ��LI�,���c�%Z��jw�+�sDLU4������)���ɨ� g��s��[�*�s	�J��P�R3:�4��.n���fro�vB��~���w�����ov�6D�O�8ꀜ;��(���n����`�΀Uk#`��Ϝ��oAAA��>'k=�����F���+([+�s��lV�E֑�I9�#��]u��E	��z4^L��4
��xe�p�-��Ӓ�ɶq���}=��1�]��AO�^��ˤ��N�?��9��oqU���C��mGӳ��F�oҠ��~�v�m��~u0�"���6�e�kk��g��0���Y��������4��o�����W�3�����a:���c��+����"0�� �<���PGr-%	�b#!'�L ���jTf/�{+e\=�eM�xc� ��(DF7�8c����<���j���+T�F��T�H9��3"}���4����;�b�VZ��^bX��Ķ��e^��<������/	�Gt��w.�ܔ(p�=�b�Vo���uY##�;%�)0��7s��zH�{�e��G��o?8箭?5�(c@E��A��<a4�8K)�H��*8+��|�(6���A��O%�Tz���`��88J��� ���ٽ��f�;�aட��-f�W#��/K,���ۗ�Tн�Il4TUt�[�fA���������]k;�J.��|��҆�O:Wc��3�V<��YdG�P9c!��S��y��~)��_o�s��X"m��DX�����y?6�\a���9Xl����V����#�������/2����͖qt�D;�씶��Hwj��u,�wC.�5�a��)�#�G��Qz�G�kx^z��� �x�7�F�Vo��k�S���2D$�l&�)�|-,���<$O.VZS���[Ldd�E&�%z�yle��N�VY[pp����l�vn����'@���U �E+�g�g�	=����~�����2���uʜ�|�����p���[I�ӏ�P����Z��������������+���BB)XP���[�LӼ	bY����>AǠ�q���ٶ�tC���gtH;�4I�ם�
�x�$h)��ﾇu��bگv�v;|� -ظ|��.�h�@|.�Q10��bn�Z�Z��?�c)��������K�:&���|>�ʂ��Z��V	�Kȏp~�MD���8�`��4�ɰ�5�(��(�4J�����;Pm�`ab�8���� *ޔ?�b`S��_�2_�PC�Z�|d��L��\��n���1f67�D)�Z
�d��)�&���1,�j���~�{)��ݕ�n��m�69�I`JpʽF9ȷ��j2���]r���������~5�3�y��օ�w�C�T�������������߭�Z<O@�14���ŎK���G˭�� ӷª� 2v&��̽��\n	�����!��΂���F��ohWm���WDf2-�5���J9����,�U��z1�B�:����B�H����b���U�/�g�xq��S��-���9ү�,��_l��V�@�w�
����|�������ih��U���4T�ȁ��r�k�� j��!�G�R@6_]brbU3m�=`�&�i<>2����?��}%/<���zg0%]P�l~VC��W�ygT�iX�X���d4
�����w�)�����6%�����{ǯ�EEk�"�#�2%�� m<渥�����0�ס�7fv�d�#t/o٭di�@���j��x[BЛ�HX�>{���ܜ~\V�JB�O����4��cφ���;�o�@ϲ����q�d�'�];O�O�@��x�1.��I� ��˚O;���e'wW����%:xB��n���Zmoq��(zF��Y��S��1�݃h�Y���ۏv(-,�2���]�E�)�-�ٻ�������;n������K"����hv��2���O�xE�J_0�[�����R�� ��ҵD� jYJT��ZԨ;���=Ũr��J-���`Ѽ�.m�ω��F�jl^�k�߽ڻ�gA?a�o!�VB�ǌ��!�H��ĝ���RR�V���X�!�	>K�["�1ʋ�����Lʌ�)�v���c&PA�3�?m$8]��Ƌ��	�G����O���0���߼����T��~��P4�?����� L�����;?X��
\���,��1���2���r�l��_�,��2aFFγ���8�y#!1���R@��|��84�?�G1����2$O����1�oyW�c��Y*�q�����\ �Q�ְC��F���?#-����#.�ia�K�31VC�(MPi�
����d~�;��>�
j�f� ��VW�!�>����iVJ���EL����{� s�������ׄ����f]�tu�wɼ���2��C�L�%_��������{:���~X�l��

��8<#|#<�O`D�z����9n�� F��yN����`}������' B!�'�5�Z���x����-����+�𓮷YK߇��T��8\j�.�R�m�G���Q�fI�h��7�ڶָ�Ju�.��wr�q�E��>�f���P�;n�R'b�t��q�T1�n�M�S���D��x���W|s��(�ȅi���!�n�5쒨ק��T�XW!��٫�_Sb>��ד}6<�q��џc�ꃘ�t�y��
�,p�4�t�,{��X����A��-H�8e>X���?���%fߢ��F���3��y��7�WPFj���/��CR��� �����MF.۾�F�)��p����F����0��c^=K�����0��1�Y9��ǉ�sq�����]�׌�V(���|���?��cV�
]��}[�A��³�����5�9/}
+�O���J�0�
T�%��%����<΅��'�n�U��'��Y;Ѝi��vv	%���qZZ��*'��m6�6��»���&��&�^��OD=���^�=t�ѽ���ꋡ���.թn�:ϕ 8lG�׬/�C������N�liS�WM/��4�[-�ڲ2������=�$�'gozz'}��f����X���<w)/�$H�(�q1���맘)��X!�$�I����sh��g�b
'�*)��ɯ$b+nŎ�Do�z#]A�^Me,��Pf٩��sP����O�^�$�-P��,�b��p%EVZ�%3������%��]|�P��9�)\���"���g�sUz'��Ǜ�TD��#�X��,i�=����$' `��4��~_���;����'���o�)�p��=�Ju�Gכꦽ�L���QJ�t��Ϻ�W�T[$}�h��:\bG���fg�/Fy?��c�q��Լ"�bl�`���="�����ݟ/�E�Վ���>����=!��ާ8m�U��X��Qc����]���b�G�]�6la�|���9l�@h�
�N=�T8�Ά��Xs`n4s4�����Y��<�s�!��by ��
/}l�8s�t���������ꟼ��s���hW�ĲUs5,F��4���x 
N.S��g�߭ ��/��Ѭr���%F�َR9h���
�4�1��^&�h�rvz����
z3tio7���s�}��o��L�n�b^R�A�ύ��}Ej��}��d�_�^?b�����i���.[#j�ڲK5CCJǗ�d/�Č\%]\\^@�HI5���q�q��-�_8΅t�R�(3@h�f)v%�At��j�;�ff�I�}�,�K'Ng�sTW$�����&z����us��~t������O�Vp�[j�tH<��󱛛��_yr�%%��}==��MM_@�m;E��vvl�������t��	hk�_!w�-��l��'�QL)�	"L�R�Z���MܫTP�7�I�R��&@�hȲ�/s�(0��B�����n����������	200((R��������𰼩���O'��<<r�Ԇ�B��d�^}(o~XÙ�s$�tE�C'V���2с�6�#i��LC�	��T��
�� )��R]M'***��5@f|���4ʍ;�Y�r{y$��V'MwU���$]��#h���P��V,pyn(د�w	2�?Hߢ��q	�8��K!���M��Y�S�]ᘬ�dy��n28�ʲ��`2Nx�g��`����{�S��w�PQQ�>1!	�7�y�=	��'����#�q�_��L�L�@,���g�y��ns�~y�{�"/D�Ɖu9sĶ�(��G�1H�٤��V,g|�rŰ�>Wj��N����|N"����qEy�d�ve�w���8ǣr�P���|�[�$:��%�.2�:^��Ja�+Ǩ���OhiG���E��*(�22(��W�/}:��&� s�k=`rQwvrn���< ҹ<ۅ�ıeK���3��<�@��-�D�OP�����C�wu>��G���V�-V_�����j�}�N��33� :!Gj�#�?�/[���/{{{�y^.E�"F�EH)�ϻ/�^�1�4z֯��y�)8���"�h]<����DoR'N�Αp����Y�J���{yb�$��XRR���#y��8m�jh�JW����OD.��.L&�t�Ugr�i�#ț����:�r�_�v�lӏ�=��4�]��Y�?��vZ6�f���.�<� �ll?Á&�g��o�vC�}�����eQa�eoϧ���`�����غ��@@��y�^Ӯ \����V�F��9S�Ϟ~�'0���wH�p�	܅W��;522�D�
u������e���u�V\z��'8)���Թ=&��:5%/����/n𣥦!�%XT��x��*�ۙ��ƧME�x��$�"�;5����ki>o��:��������*�fڟU/�����t�����bnַ���e�8!A4�+�DX�
11K� bWr����&sf��$���#���H�~����YK[������O���VR�4O_����h#9��@z�#��B�]Pȡo�9�%��1ڵEq��o�^_H��DQـ�镌������y�(|�Ή�$n�4=��G���}![W�yG44K��'�H�0"ɔ��anv��h����*�I2������ܒW��� ��1+�b|��ݷ��o$���)�[O��%T�C��R��p����Po��B�����_=�T�#ݕ�x����]�T�M�����r�s���������H����V�c]_k0_�(��6��*���Ś2�o ���!^'��$���u%�ώ%�Yv6�h��������r��ݴ~�n �m��̫��*
WW��	6����9��N��C�O%�s-a�K�z�@�4�����W�=JB
L`��Rs�Q"����A�_�8�>c2Ȳ�4�"�����0��o���`:;��M��p;����[��LXJx]i��q^!GL)�Z�g/b؊����;'A[���F�La�bH���4�<�jY]���I'�V���߉o9���d�(�Ty;OeI���g����8k�l���̿�~��?�� ����b����_S����\��b�6؈gGfX )��r�gB^G_m��S'�2}�K �4����}�[�����'l� <�D͑B{D�?&Əe�'�V5�%��-A���:��ʅ��K���(D��Df�J���2ٞ-�D�5o F�������9?/�ٓ5��#�P� �!r9�-���ڣ��1X�I"T�I���[�2[b����0�l��U��Ɩn6N����S��F�U
�/p��?_@k�QMZ�kS,V��5k�đ����c���;U`���,(����T���Si�}����p=�o��!��Ox�u~����]y?�R���/�>D�UN�"v��Cb22���>%��z�(]`��Hg9��4$z����d���yiZ���v輆3�s�#�䜄����gXM&rkA�,0x��_��cR�9����Y��u�@��<�)��>���EB��c8n#Xde��� �4H���1���̐�eDe��K��8_�c��nҚ0��ʕҰю����W�;=��kX�с)�Ұ��`��,Sx�:�ƞ�'=�o:��o
����h�G��>��z�">_��^P���>B��_��N��'���?���o��Rt��o��j�Lë�L4�憒�Rry/ﭓY�%��\��u�.]����%�V_/\���ཤ��]_4�qMi
X)����B���
�W^�7]�,'���3o�I���Eݪ�l�CBp�ա�M��e�݌����Qz��=w��d���b@u�La�55!�o��FK������ip5\9J�� R��?�q�s�X���{"�F�h�Տ�~���i�Ǆc�}� 㪨����^U�"�O�	��|��yU5��4t��ce��M>�!l�R�� ҲM_@��kB|�ic)�lH	�M1�|�#��:q}���v��p�H�s�e��ߺT���BÍ���Œ@�%��Mai��p�J,��m�ِ3�W��ۓ�-��G�{�(fp��ͱ�M��cؐ_��`}q��.e�>�\��q�����q��.�ީ�) ��K�t����ˊ�oeH��Z�S���H�S�t�6d�Y��k���{1���&�_3�_���+~4��l9��o{,�s�-��a��+��W���yix��!/{���`��{8��yr��~����8,oED!��S/�v^n�8C���sz���%�_�Ѫ#�$6�l)����	��Z��,#�'�9�
�D��qσ�Q�^�7z���Ȝ�R|EE�T)���X=<P<��ӑ���]���rG�Cc�+s�!��¹�����(d
�)@�������R��Uj��RL��>�=M'\Nfs( 	��R/f�G���#�Z�e� �����g[2��H�����Lb�W�]9���o$5��3��qo,�zh4��8/�
��v���V�� �t&�Ư2�Ծ�wa 0Cʨ�x�^(C355�_�<��+���e_4�W��թ5k�����^����[�P�e5V��6Z=Q��\w�G��bd�ߔL�m��S�D���H�������}��)ޡ������W�R����R�N���I���(;Q��{������R�q3:�ۃ��+����yUɥ|� ��+\�g�������4Z'��o'`���uK���z��j�TU�5j�AТq1��f�L���EA��\�W�
|SA_t�I 8�BQ�$)�O���t(*��3��u��ᷥ����
˘�����s�[9q��iq_��>.���w�i�ݿ�FN5�,N;C�5��F$�ewe.=v����k��o��ܛO����Z�n2|z�q$\"�#�ʑ��5+�Eo��%7%{��t�i�q�a;�v����R����:�tI*>Ml���<��q�MݖF lt�Yȳ��h�����v���	K�%n���������K/6���Zh�������>�-i�E휟�5�NO�t��%�3�O������vt�tԏ��Uf��/2`uX��԰�0.xp��͖��2�Y��R7��t���Ł�Z�S����xM���L'vG��P��ox���#Q�N��,��ߍ|���)�t<�RX�A�Y���M���7��MZ|r�+����!����.?=@��Pf�UK�v�|Cb�!y����h���j�ꤏ.W��$�6��"�cï�T0�۳0|�����kȘ\�2�	T��(J��i�v����w�`���t�����<V���w	t��'�߬�vj��=v� ����>G����7�yh� ʸ��Sū�G���M�T_b�'F9h����Ȥd;-��V�!C�y�k�`�iew夛�2��`ʎD�����O���Կ�ZhP�Q�;XP�]�6��1�  ����8�h4-gմɍpl)趾��?��yC���7�h"�Qeۍ®������*"G��S��X�8�J	<2^Ù�G�8�s�S�]:廧xq�]���P�!��g����,U�5	��l��q �iU�l��z?�[��<���^�ql��3�Y��n�"�1�*�<�:t��
��eG���)����I:�5V]�%ù»4C3�]�+J�!�l�:IgD̙
kB]o��p-�ㆨ�C�ɟ��'��j�c3�q	�g�P�rEC5��h0�ق/���H}E>Dw^jaB�|�(�=4����G2+,=��S2IE��7b�2��y�sv�hu.
P�	��w}]�jh�K��2J�^W7�7|sC��>r���܆R$ ��év��#�&6�?@�(���p�iu���!�g��<s7����7�tɯI��N˛a�`'�+���"i�z��xXw�{[���OE��u�<g�kwOH�ώ(�:M���lV�Kr'[����[k��mdS!�c��L(�/V8o���q�9l�Vʥ֎H`@Y����ʺ˘&�I\ ���������(Cmp���Rv�o�7�r�Z�n7�i����4ު��)��\p�:��a�� X dU(Wd��`�IC\_�CS]�D5���P/
�0�е�S3���{�A�>$�뙕X~!_{���d���D��ȘjEc�%�ދ1R7��e'��k3���4����Qx�W�1���P�z�#s$��Kw\����4���!���g��+?����:�ܑ�7�[o���.{�3ȓ��7�� ��&�:��&h7�����)^�x�w)V,8�Ж�N��]�MKq�[���.������ߜ3;;���<�s�٥�xHVU�uj>�	��{z�C�UW��h���$���w�\�i�m�������:`5u���)���L��1�3�j���_��g*C���ݢ�l�V= �o���Jnj���`>OR�o�-)n	
j_��ޥ�r`���OS�]�Icd�e�+��Q��� � ��`�TJM�t�u,��Ȗs���YlOg���Da����(��#����r�M5�[v7,���M�_o�3�[�*��-���8���Z&Յ?x�vb�w�L0܆ ߼�B�����q�@nW��N�n�;d_�F+_l��/� ����D��ݲ��B�tZ�6s�I��7���I�H,��W=������0�Ҷ��D�=f����1-?��G�Ș����w�MJ��)u�� ��lH}:�/|�0Gr�4e��|k�U�I�Y�6��h�aC|�wB����� K�/]\� >��P�R���`M����4y}U�MC��6���Ns�<�տ7C�p��n/Gg�B2-�.������
��ُ(����#y�@�j�.�R�?'f��;i��&S����c^�l/��2Na�\���f���Z��u��CD�W��n��	G��Xe�߆U;b�1>oe�%7�&#�}&.���-i���]E@K#��PϤab�쥌�����pO�*��+0
�qX_��ܬ�9��,�i�l��a�M�gh���і�J��B�Ue���4_q���.N󅓈��;���c-��t �|B(����P??%姞����%:�p�����W��z��E*"$�x*��e8z���w3zZ5Lnk.f�h�t���H4��ݙ�kr�1W��Z���[��ȫ��i�����X�a���Uꀑ���N#x���|w�0w�ɹ��B{���M����ѐC�/�ʐ�� .�4 �����f!?Z\I��E������Y�lZ�A��U��J3�C1Ku)Z���kX�\(����;f{�Q�oM��(Z�P�-�6��b��F1I���M}�k�g�qvI^��(WPm��=)��jq�{C�uK��L6�/�cWEf�hq5~��hI�'=*�4A�2ǶsZ+#������QD���G������?�i�U���g^���8�֞�����"�= y><���Ξ@����{�;��];ЇY��i�Vu�#?�\�.����6�T*��L���+����1Q�W��m�v���4&�)�a���D8|��c?�t���?�El�d5�**H����A�|^���ğ'n���]�[��#�K&�Y��	��ٕ�6f���j�]*U�]���������b���u�_����$�k�a*c�F�\7��7_ֱ�����O>����T�����	�Έ�l�;�Ph=x�o8�����/�⏙������b�A��9uJE����$����eY��4��7�w/,M��BC����<;	 yjYF��[.�-�����0�*�����Oۇϛ ߾�4�|�ӛ��T��G��U��O���M��E�i���M�~@?f��4���N1�MQr S�v�ڬC�r����x0��Rq���gRO� ��ׄ����HP~T����=�����eH��I:bs] ���i^��V��T;��ϻ�*��}(5M%w�]�aX[�5�n�����S�k�n|�)NJ��%�bʀ����/�"���7�$z����đ�Rz��a	Ξ��.J�­J F������Y��]�-$=Ν�����:΋�ɷ�������6�b���O΂Yi�9��S��<����`"Y�^1��-�T7^�Q�/7?Z�}�C&���^Č�3|�����BQzѻ-!��'ا��G����l�$
�(6sH �
��[g6�s����ɡ��'笙��Z��M�%+/�5�(.��	� �Z4�����x�31�F8B\^�?���DDDj��?�	
~OL�{w}������&���E#�K`eeeqwu�wo7[?Ń��Cg��3b���N�o��u����9*�M����]��Cu�DX���XQ9�����;)�d4M*�d��JD�����$�\�r����3��:8`��̋�Beł$ �$y-f���L!��W�Gҁ7Х6��ҹ7�l��!�W�+����e�:�p)�����y	��|����2@peH&ǧ.�����U����Q��?W�?4��NUL���=�熭�r��W9>���[�֖b��;lu�\��f\5>�H<���_6���\��O.~�}]�'�'�����M�a��Y��tG����K<�%��M�v��o����bCE�Ϧ���	�����B��s�o}�"l,b���!HW��Б<:� �ǻS|�&RRRJJ������J�]��冤$���7��}GV�nq�̻��F�C��1�"�2ŷuϳ#Q@�}��H�rwN.�F�f�	d��%�i�c��A��] ��~�	&9�I��t�)g�Z9/��`���+��W�W�l��å��E�4^�����2/3��h�RG�K�j�\2��͞	��nY���xsFd�Ǥ�Ȣ���$���>�m4��������c������M:^�.,�]<�Uw�'��૫'~�R?�Lh�b;��Kf%q�S�����?Z�[��}-��|o��������fn�~R��������e���A0S��P��.׫�u�0�/y|���]�V��7�	e�CɏX�B�/�p"����&��^�ä��s)$��aQOg8y�X_��8�tfl}�+�V��'��?S@�
�-�1Y�:/ �Z���M�q3���yr��m	J�0L���D]Gٱ��?�l���WK��������~6�T�HD�6���8��"'�����^��*vR�En�6p?��e�������_a�A��3͝�]<�t�'�c��w�LNk�ݙdB���gm���:��;U��__����>s�<���r۽Ei�e}RfQ���X�ܧ�A��l�K'2dO�	�� �Mp}��d��w��X��*��j�\��nol���UXUX�¤T�epP��c��������<�����27ǋ�j��֊��n$X�L8WϹ���Ԭ�w�>
��7݀W���BU��f���&)ا����4Pq��������G����7Ç�1�@��6(��+���*#����p2�	G������R��ͩ(��"��I?�l��}8p��c��B�%[��ɕSΕ݌�F-�Fȉ�s�Ś�Y�Ǵr����"�S��l��R�k��K�5�D��ո���Mm0)�^��6E��߿
o�ؐ����Jy.����v�e�˨��8OOO�c�P}WG-�pP��J�}�Ù#;��Eჱ�!��sb8�ծ�-c��؜w�k��O�/P~Et�;k�j<A�w$�t�/&�V%�*�2Aw?�f� �)�K}ǣW`�W�0���0�p�ծ���1�"[�~�9JUU��ѝ����6��JcV�β���s�8����BgoB�����<�X^F�J�F�i �p�Pӎ�hb"�q�~�~ :[�n����Mz�ҟ��=p���蟢`��������>����7l(d=F�=3UWo���(H�~��o�;���l�7�j����^��8��vlFA����t)J���ꠘ\%�u*"'�*?:1���@���7{L�k��D8�(��|]yydTK��ꇗ7�Ǯg*߃i���n�쨼�X��
���zZ**1��7�c�y�?3d���F_m��w����8O����ز�4$(���f���)|�c�9�*�4�V%�ߐ��舆\���PhZM�tnnn-Sӷob��6�=���;;s9H��{������������1n�k�HsP���,�L��Wx]�Cz��!��t��Š�	���
�/)�hzx&�(�����/��YYY�#J_�+��?�!��÷/��P�nz�
Io{\��{p���R��Wh����-�C�4�7a�/N��f�m]�����M�<������~`Ց 
9�?�^,���� 
#��Z�g�M�F��=�Cb)�!{e����� ��H�K�1�a�����:y�t|Vir�'0$P"�!��	�E���!�DX[%�Qm��#]���l���o�\��	�Ì��p��80��M�<�l�,/OS�QT�~���grk�(R携$�'�7̠x�X�R�W��2��� w(�v��T��ݺY9��X�&�;^VJ����xʝ�Z�: �մ�!�U!j���>
@b�'�E�jp/�u#Z��v��<6�$��^T�Q�vG;��W���E�C�@ �K)��8��i��х�f6���3�����J#c��{�n���HA�ór���)9�U1X�h�G�}��F3[�,M�aIY2���[ng���r�nt�)�R\�g�P]S�b8�H���"��Y�'`,U��RG ���`�z�v�[m1����
��x*�6D�#-��[�X*^����_e
�����{�E2 H$N��=(B�^�z�~B㯧�'Nh>�ǲ�1���o�
Dr[�1�2���}�:?b�5{����1y�j���ВT!=����m�Nڹ�o9��NX�wr��C�ɟ5�K٭h�+X�5�e�=��G�.j,�~D�%2�m]��<Pu�N�@ʿ�?3�:�P TxNayZt[��<�פ�`.֪�q���y��Ɉ�Zu�<&�����Ub�0 ��;��ՙW�C=5���6~od~�*¿�-�����әB7{�r#�5|��}0��/�-��ѥW܄�t��;��=Q�f�\�K�f�����S�i.�D>��LM�T0Q�f!��5�)�d���;y�.�-`�jX�_Y��9�wN"��\m�ұ�\�����ʽuWѾ�p;u�]�L�i���	kz��+$5���B� 5b��u�Pa1�K/1"/D� �2�������çTo���vOxNa���R��D�e����z�ng^�T�����W1����M1�E��#EluD!��y["l��X��2��� �3S窼Y$����r)�E���yHC�������<�N��ޖ�XͽXDZ���(���/]�����4�|�ӹ���}������ �<���1Yx�P)Vg9��گ�-�V������"Ү�~f.掊�e�������?��� Af�p��pi�ᔒ|�ک���Syz��`��s��Yl�P�����ʶ�:����9�����a�H8d��gϗͥl�oG��� {�]�$%�vJ��l�FE��fl�]{�&�PM�k�1'm߸W�Rt�|�rw9e��Z�'�B���[���	���xRc� *2m�8���v��dRb��fpȣ�����f���ʙ�|TH?̑�Y|��@��I���+ݤI�}������f&��hkhbh��p�?p 6���yH�b��մ>Cї�,er��V���d���z�[����2�X)N������r��I�vBRI���^�K�lBhf����3���n���"��wܱm6�o)���f��P/�I���7�Zl�a�E\3 ��rs�&��T�%�/�X�S��:�'����onˋz<�i5�Y����PM��q(����\2���9��cϹ��{�����H�(�4zȻ��?M}��[�e���������ƴq�t��vu~/���CmR�w���s����M7����5�yo�g��Ŷ��1l���*y�$=�$���l�U�PY�Ey����W���rĔ�q��kj0/.'������:b~[�%V9�B�7���6G�-�r$�N�Z�z{�b�t��սj�,�j��6�{ ����q�l#�-i�G��3|�-L��c�Ꮢ�4� ����9�Cs���>�_�U|o��T�_�F�^q��Lz�h�Q3>_�\/�ɽ��WX�1�}U�	m���w�Am09ɬZ+H���ES �s�P�F��?��`:�#~o�߬%�~����6�>N�@�3Z��xWӈ�6�lՅ�5E��H�Ġ.�>�T%�-Y��3�9�R�������XN3 ����0j�E�/|u�8|bf9ī���x�p��]V:��c2_��9���w
bކ>g"�P�g�H�zX��������P�/]���WH. JZq0;l��5�ReH���&�&��ݗ��}O#c�ͺ�����E�4�����O�f��I��dU3��Q��Y�����5�?��`�_���yv�)Ł���oA$i��0w�����w@B��A�p.�;hj�s�vl�M:���]��wB���sL_��b8��~� �|b.�W�z �~�R�y��L4�2�W��fp�t�`!�J>�����h�[,����7�[�	�<EiG�6a%7�:FJ5���r�=s��_g�o�T{[x���'��Q���qȝB&�o�Ų���`��z/�8��;=ץ��L����i�0n��M�{k��Ա`�E��j>r�7�	�_`�ÚN�\��q�b<hm�����O�E=����v�N�B�d����ڐs�e�Q�[aʴE�DB���E����5��<�8jSy�k�b~ҵ`�Ԝ��$/�?V@X;��W�s
��}��� $�O�Ց���v�m����U�biz[-U���;�&�����:[tw��C��l�����'j��Ix�h�+�X�J�1�2уP[�fxmX��Gw��o�0B�ozn��D[/B�Cl�+G��j	�5�pl��^��������j���h��폗�����g؎7aY�D�,��7T���I�����S9�,�8�l�����E���o��9XN1.{�}�z�E�	�)r�,���ѫ�%3��S�R=�	��?�~�܎���B��L�\l҉��;��;'�sr�?x.N��,��>(��{��E�l-�%�)����^��O�Ǧ��d;�_�V�/��!�7�-��R�@}�]�{�}	��/�]yW�xH���N���{އ����(����������
�ɮ�8�j�����*fQ�y�������I�>��L�./1m�6�B��٧��I��,3mu�J�tޜ�鯫�nn�vqa�ǵ�i�a��1�kH�uWȊ�3nb��ȫ#Vo,u�oRan|�y��
��[#��D����$i�u iE��5&]t1��U�y4��<)42����~�//����W]���>u���H,����D.���$@�K��E��C�*�U��^��k�{��"��]��K�<^iњ3��_[��u %�l�<������������g���a�
e^�������x.���V�(p1�N�4Ê-uS��f���/�����}��-<>"�{]��.u�ܶ��̘����-����,dPN��0r0b�Dc�.��Z���!!�=�3�k����᫺@�F���鼰�׌d�e?:W����p�=�>U	ݮ��|UZ����S�r#�s�T4P�k�ltȸ���S����NWP�ݝ�"\���<�\	����T:�O3Q)Z���g 3��g���5� �F����0q#�����b�B�O�{=�嵐����M�z�F_���/�����I��^{Y��q�/�Z���������J~('���R���Sdp���׾J��q�~*O�0�Od�U�4۩G6^yi���5�c�*���
om�v��&��~iZ��Eߪ�q�$��_@����J�[7�����m�*��1��!㏦�=
L�X�kҡ���i�\��A!eˢ	��D�~ ������ �gH%�Yժ��,~~��Bs��08��<Ь�ڭ���2�"��Ǯ����[���mE��{kr�3U^K/�'�����]3�G�3❳T�͡��f�v=?�J��m���H4�z���)R�تq_3�߸�RB���ڰ�����A��m����<$�v��,����	zt�qzd���&�e���O{���%���0%��M�Ⱥ�ՠDg�-(�8fI�7Kܺ'I�x`.�?���li{�H��r3�*�Z8�cC�/�
���F��7�v�s�g�H�C���ǕT-3������6����r����8�s�lז���h0��Iv����۷��w�V�-h��X4l�e���mG^�h9Y!�,��O�}��>NʲA\s�Xg��6g�
��w�c�,NԿc��X����� ��E��8Cr�v��ւ�'m��h��3�f��,0�l�L�]��#Vv��M�A<��e�Z����ؐ��˫T|8
�5b'٬��J�7S��e��o!Օ\�t[�0�+�јed����şE]J�Tq(3�@���@�ECS�h	�C*O�tGD ���� �{	Q_:�G��_�^5� ��a#doA�!���,�f���+>/A�UE�#�
Z��,#������ �1��K��M�Q+��Q.As|/�%�R�J#s�WoC�H^#A�������'�"PQ���I��p"� ��no��r����Ă�;%�/���,�E�gxR1�/���1w�i�����[��%���_�{�yKWK��?N�x?e��~)X@��x��[~��.仳U�/k� h��ee����D��w�'u�� $ Y��p���	@*�)��[8֕��2�Z6\E�g��bL$3���x��o�3F ~��%AiT��r�)*#cx�<D}� H���Ӫ���dS F@C�j��?Ic5�8&@z���'�a�&˟��ED*��Psgb��K�P3� �4:'��l8����Ϲ!g���/��"��An��3�����?K{��l?0��̋��z�tX#��A���O����Z5���	E?��11�鸝Ey��`��g1:��6�0ג3ڝ�^T�Tu�h��Y���Hw�!|�eZ*�8�������Q���������C�0�6ʭ;�H��H�j�*@z��>�H�DnO�ʣ���{��$��N/`�8]�%�׮��l�w/2A��
fŀ� 9k��+�vp�_#T�� /9o�~IH`=�zc��yM���Q�ğ�Q�|�<���/O�s�FH��i�0��R�F���V�W�("���"����R ��O�-��}��V��OZ`�?�����R~'"��4��܆1��߿v�+"��5[(���y��H��pٍZ\6�[��U�ȜcQG�0</!�x�	���2��p���Jf��}O�3�FG�U;k��b������Yl��	�?�~6ϯy���	���7g�l�9J]n'Q����x���_�k>��K$?�y���;^v�n�{ɑ�J���峲%//C�����V�N\�L}�����ۚ-����[,�W�������~��K�-��F�y"0�A�';��!�VU�H:Q[�O�k�SWV���DgA��
�y����s8��߉!��m�Pf�<��M���}2������a������So��%URE��a9{K��/~٠_V���o�E-&�?�2�a�{fU<m�[fh�溛"wC���*Z|�Q�m?r�\M��c/Sǰ8�]
�浺�ɷ��9}�*�L���#v���Z�z5���<45G97G=��`�w����C� 6��}_k�s�?�b��m޲�����K�a7�Ca�f�{_X�(�u�Yo���a�I�;�x����Wa��a2�7e�� �c�!0�����������s0t�V�Xr1�)��ÄA��1��7Y��I�H8mo��ǒ��L[������u�Z?`yܳA.�C�p�����^:9�PY��6̤��?z�M�k���1�eB�	�P&��P�8Y�<XL�m��\�_�B)n0c,��NŰ�u�}a~���,�X����!>fCc���L���]K��f��'���aRVNXp����v�W��թ����2}��a�u��P���j(���o�U�f�8�9���$��-��*�)�_���ヶ�ﺃ�	[�q}����Z����Ѣϸ.�S�^�kJ>mNM�v�Hv����n�j���Qj-��7��<TR��i��@�]��a-�W/��[�	�5�4�+��=��DΛͺ����bQ7
�.PD�8�rƪIFT!���6]�}-.���M7)i�s[o�}<���ü���D$����	m�6����@�cmQ��q���u��%�GG#
��gQ�j���[�S��Q�d�Gpo��~sn�_3�l�� �=��ʣ��;8Z��+&}��g$��SXq���@��������]k�Vz�$���U�;�)&P��$H�<��F9���`��x���$R�4(�c{�p(`!�4R( 1�ǖ�}6q�?�D���2."���MA+��62q/�<��fV���(�2g���& ��D!�ro^�e��xV_�t	!��8S��qWqkz�EB��D����F�K!{�L�U�]���GUt��z�ߥ�1���c��C���ȫ���t��0��u��=&|D4$���ǚ�(6p~�|}?;�1d浚�x��i����1&.���v�06@��Z:����
���/�ƣ��8t��@(�Y���g���O�a�Tt�`�W�G�%S4q�Q�.��5���L��A�`X���_X�=���еq��~�L+ִCgX��5aV#>�sFG����>`�֔����
4�b��"�·AQ�WcB��ݜ�E��s��Da-H�o���w�cT�2^�d^��(��<���lòj>T����#P�%���+#q���A9�9o*K��A�V��RK�>����\Ca%�����k�j��f+�#��m[�w2�x����J�$�P�j@fݾ��,&�c��d�K�T��қ�y�M��_PnN�l/�E�uu�o�n5��g��1���m�`pΏOE�� e����r�x�u��L'�G����}�X��'Z���Y�hcm[�Β�5P��E��Q�pw]�E�E'c܋e��;ЊՊF��g�L�6*f�W�3Kh=��jY�J�O>�����G%��kӣ'�+|����T}m_j;2#��O?J���ߐ<�:9}mZ�;Md7�OB=6�>��m����Tp.N���7|AU�J1]B
(���5�P�Bk���kGeɟvN2M��R���M|�Q��)�9�g݈��.�o[؃iz�wl�ar���_̑sCߥ�����;��|�D����:K�����"4�
v�}as��@��6��{L=}1!(����$I����G�Ja���m� !��+3(AD@&���I;�k���{TtM�>$���P�=lB�]���S�U�7��=�k�"�.��� ��g�+�1'��������&ν0�Ԇ��Ə�����Yc��BG�V|J�M��&?ʥ!�z7=&N�&�~�#@�=<�ɳH^>c���j~4Z���X�e��Xo�3���ڼ��p���S	=�����6Ɔ��z=4�^�!��;t03�k7�V#�0��&�/����)���X�+vB>+�z�w�Pm&�y�J���x��.�QdW���J���6�FPR�h T���&���j�U���N��O{��YR���9c��Q��nExV ����~���`�S3p��		>{\b6���7��F�5�dk�O�O�\~�QIA��+@p�5Ɛ����,�b��G�t��ؙ>�GW��������}%���<�]���^G���^%�8�]{dH���#ڧ:a�N��UFqb��\\u��a��%��#��L���C��)ST�\�F�W�]��Sp��g�M�= I�	�P��;?��*�7:����W�+~׾xa�a&��?�-�Jx�X�$��� %/�0�F��o��?_��<rZ�$��}����:�I$ADĊO������Yq(�����0��^]w�L#(wv�t�rѷ%�ٴ'YG��s����ϻ;���_A欞,s�7��ln�W4�w��&��S#�/��@ǌ�Ir��_�d���~巙�W�a�&�r�f��^�xF����$*�*��{֕&�ɥo���$��	�l-�!�/�`Ҝ[�Y(���IS����&-�������O�l��Ou��'v�÷��c���j ����(��#����y襜�dփNPFr�Bu�~�,��"����_�=��?+͇�M�*��!���6� �)1酶�@����[0�w����V�:�L����͍���������x	��*�8��w3W���w#�*�:���s�W1^��^��k��`�X�I�����g!EO�J����Z_�KJNP?��?�:�>`�߇� ����"�IƷ����Xe)��h�����ev�~M����}��Ԝ����y+�&�HG�jE�^�nH]y�,Jd��� �����c��~�t�@@��̇j��e_�<���yD�����}t�֑�)�<��P'F�$����)�Ǟ9��z����OxJ����|+�G��(5$?dj��W�8�V .e���3#����)��K*}�f�~G %�;tRu�AW#S�n�;k��v��%��.���%GsRξ�s��	qMi�U�@��l�G�?���R��%�۲���мW��:��.Ţ�?:��j�r��ӳ�����ϲ ���˴¯Ǽ�m۾�*A9���$�@���4� �(Ԥ���}���vB�zBh�&������T@�p/��ډ�R�ק��T4׮��~�;�'�]�9��e-��A�T��5�WW�����sA��r��x�8����s AE3��b��<���2�Z*�����퍒R�x���oz�, ��<��̺���5�;2���Y�U������ ���C���4Tr������7���u���D���W�ªҊ
��sݸ[߹:��VNA܁�}��`���E�~B{=��ob4�LC���3����nnfCk�J��g4룞Y���׫o��]w'qo�O��_���؃�.ݚ8�ߥ�����\}O�&
��@�"ϙ%y�H,Ю}J���{�y��_��Z�9 �A	���}�
A��<j����0z��cM�{��7�Zf���ZI�_���Ԃ����IE@BF��������A��hw�#G��c�_{��E�e/�}k������g%�4��&��Aru��	�\��p���S�bs���&p��/����d�Vp�{W�'�'�� J{�Ӳ%�����KJ��Y�C�ȓ�-ׯ�|!	�8XX�7�]��xh�U����乤w8Kt3�<�~jx��Vx۫��޷0��`bbR�� Y,�Z?Ӑ�(����b:u�A/+3�"佹�Z-�����$�)6�n�$�&�T��}�e��[�m��y��������%��$�i;�,�3��I\HH���v|tE�rXjm�E^~��4;k0�,��t8$.(�||��R[^�����ˁ2�'q�H�KAwo{�9~dEi-p${�\��$��cdnn��=�6�
���CCQJ��$ֿ�f.�>]=^�}��xs>)�Xk�0�#���0<n�·/�G�xl��WUW����͆�Xf���ڈ�9$p�u/W�*�ܙ���#{5~r9����،ߌ�10��v�B�Ҩ?e��U3��Zt�����r����z�i���/8��I�!?���o� Lt��%҆ml|H=�IT�i����m���;��L��#Z�QW��㛿�n!,B�$��y�9��J/�#q�ю:.�}����1\;�S� w��+x� 2���O=C��=N����:����Z�����(�|�٢6J��`��P70��'X��fg��3}k�2Vg��D�qr%����"���s�ԶE4�Mj����+�/��q$W�||��������L�,���?i�ҽ��҇K�#��0��^x��*w5��'���c��oR�8M�G�����ut6<�F�ٿ ���P|R��oVu�=hv{ItRVuF��	�c�^��B�/���LMiO��x��~$X���+����e<�C�'o�����]}�WF��6��]>@�O�D^�IL.����U�W{�(��Q���.ͮ����D��|�"�Z��}��|r�>����tfp5�oΟ�����m�D"P����'h�fzlBB��"�6O^��^<�'<��m7�5�*�2;��V�Z/㥚��i=A4]��U�y�C�c����hD�D�7l�	W|����N_�
g�]WY�6���M���z=� ���%���+�%��V�䃔f���r����q�[�������������n�`e��Ȅ3�,������U�A���M�B��b�w��|\���M��G<�h���r���!�o2!bQD�]�� �qo1���.f��a:}M���SPZh�s�,�2� �:���ǈ���	:����Fɼޞn��&m^�|��5|�I�,�Ϣ���R��O��
_"�~��Di*�i��)N�R��F .��8b�K4�+zT�'zTcv{x�F!�"��9"�]#>�^ՙ�Nss������RCsR���1�qr���rZ\���3Y���3�A�UFI$�4�6=�Zj��`<ǋ['A�Y�rH����>��Q�&d1���%�1�l���2D��q����oN�|Wri��A�%����m���iԜ�zs���7ʎ�����ǯ��<q؛���~��'w��5]�����@��� .�_���)W����UWp�U��#�H������/��QN9$�|^��Xץ9�TP�[ ����z�?�����4��m͝R��1~�.ӡG��U�~G��׋�Z~K�2��G`��C�YQ�ٲ���w��ׂ���Sr�e��/Esz��4.� '���!�k�
H��~�㟹]D�ls���T}>��H���g\z˱Y��`򛟉��/-�.���$�DgS'ފKxo6ߣ!I99p:b�����/Z`�hI	G��#
G�7,&9
�����> ��l��,ƥj*\��n��Ũ%j�=�E�:Z�]���B��Mi�R���~�q���4���Z�w�\y���P�${��ޥ��Xw��*P6����P@`�"��������G�?EQ��j���cr����@����E@R�Q"=�4�Zg�,���Ro`��i�=�ΰQۈw�^y�P����0:�z���VᤨQ��k��°qO=o�/�]����lo^��'�0jL��?��X����/��C�jӌ�z�����q1C��%y����JCĘ�e;�y�3�B�n'YQ Uk����|���_�dC02[?O�̀��ݎ뿞`��#��6��-W�8��]�� �A��i{�����L�u׌��������Ű�9t�g�.[����S%��7���sx11���  ڒ�Z�6�����kp|��P�H�"ȅ�����6jA|���c�a����O_��w2ˣ�T��K�+��'����[\ }��P��pf��;��z�?o���L����g�W�K����7LD��10�ͮxv��O����Dn�+�+�V�d��e��ߞ����K�()��Լ�"�;*6�U�#J��/�[���bIE�
�#�,�5�z��%h{9�\���fÌ*�WE��ï�#[�T��\�`�����x�/�y���q'��o_�^�c�u &�T�w�6H4)��n�>�ڎ�A��Hs��Ʃ����Ϳ+a�z~��c�E��\�@��+cZ��eM�n��5c�棉ay@�?M�&@=�]$����iŦ�Վp�=�/��F�',�xo���\5��K�����cL�Gi�waω�mGϳ�1���6���&�K�?G�~��	����͢zjN��p)%3Y?�����W���GP�^͛G�|��\!��DvP��`�#�~��$pY���C�7PVu��*��cv���=�<��pP�_��1L��Qp�0�u�cx_qE�m1���ߝ�"&5�� �:|�g�Vm�4b}%����ƪ�QZ��0���b��Z��<�R\�������[}���O�m;��(AY-}��a����33����?�SS�r��l7��>�
��p�g�ggZ���:}�D@h\�|
Z��3}*���~	aa�a3&D}Zuoj��e���;������[��s7� ��s����k�����3��q�� �J����,���qPQ�W�C�*~Y�#�9�hf*�p�/菴����|�M�ĥ-���P^����E]>�/˝B1:h�t}�O�_��_�&����X�2�HZ�����ʳ �^vw|�k(� 4��E�܂��C��Ό�0"���NuG�f��z��<y�m���`�>�OkS����DR̗�?��RƳ�J4g��R�R��`�I��F�a��9�<u�(KBI3�.w�����^�
#��.�o��$�;|�R)g���Tm��l�QO�5kŨ��j�l)j�R{���+5��h�VT;v��֎��*b�W��;�=���s����s?���������k�`���������������(�J�Q6gl��_�O��.�^��skJq�Ht!XXI�A�~B��.�o\p8_it6,�C�>�|Ěrߴno;3�O���(��s��-������'�Pc�]eϭ�6��<xFN[�l�^�JAN��B���T�3`<�����Ѓ|2k�����\2���i8��igkZ��)n�����_k0+������.iF���-������ %b�����3$H���~�4�'*E3�bP�T4/��oy�7���'Qi�C�`���DU���:zK��,)^ʷ a��5�69)m����J����([/���󭣀��d�,]�\�[J�-X�g�魬R�爭,1��0�n>���pTυ�o@�d{�!��߽��,L�v��<h%��-1���/�hY�>�KGI�Z�1[e;���1,e����$7�(;�,.�q���F�d��3��IL�)y�N��`��8^gB���LV%��s;9�e����7���N!n��y�wk�s����\_��������;qR����P11��f�b������k} +(߳%2������2����"�,4�r��H䐋��:�$i%�_b���#�HZtoR��9o�Ҵ\K/�jܰ��Ⱦ}_*z���N'�b�����9@3b�!�Y�3��%�(��3+9���i�_��2o:�j	M�8��э����I�קQb�_u�Ѣ�p��I:]�����/���ɡ�qD�97�m�!o�f>*���ޅ�؎�rh��v~T�E�[U�qU'_�\�b|ٯF����ā�z�|R�t@I.��2��!����%ފ��@��j�h�_���;�9��:�K�%H�� |�-0��� ������Iɽ�ި���<�G^����6�i6%��"��v`����4���puM�w%>�������]��Y���؃�9��ң=��O�w��INob1Z§w �jP�e�3����A	��3�w�3���&ƨ��QGR��WϿ�mZGNa���ߪY]Z��N)�_ʇ:	2ᰡ�pr� �(�9P�(4ʲC�ԏW+����,����T�˂W������g�щ��q���n�s�B*�n ��MU'�����KP֧��,�4�7����:�A3��Ru=�$���Q�����p}"P"�q��B#��������0�ɶ��w��yQ}�f ��ը��!=�
(�A�h��]�t��X�+:�g�fa[��[�Q�u�<e��~�K�>�׵��������M:Xy�-�}���{��!�_v�߽�M�G.�+�Q����<dѭ�l�WŷJ�ȃ0a���������uE��[Q)�1�>��L
@���GPcw�1f�]���h���7/jUES�S�)�-���'�tq����Ef������"�r B��'��{���.�6@�g���,�@��Ʃ�MlU9�U.S?��ua1��ʇ���G��sLX 
:��=����1�<�[��_"���&�:���ӌͪ���\���A=�b�C���7%���"�:ܔ�,]��'�K�ݎ���GKT~h�14�'J�VN�2��d�3�	^�rP������;�L�dP�p�)&Dyo�J�8�ĥ�1,��#�L��\>�^{ы�zg^қ!�"4�o�
'!�%�'�@K;'�˅����y����i���};)��3�^�_�� -����|��u�}�d��T[/~@��f�8��X`�j3�!dpAe�sqѸ����\��-l��
��8��oo-�aB���~v6k�8T���v�i� .�n���Y�e6K0���0��KF���a�F{�i��[�2�h1��X���{͛�4����ד�����i�b���1l�^�4�: `&Ȏ�7͟��Z
��ٷi��\����u��)2^C,�@3� ��ev-:�Rwb�BҦƛ�a�<lVx~�(��!y0��������@6"<n��������'#)-��cO�f3�3�����]�loC8u2B��������K���-8I&����7�kx�Ǆ��� �F��Ae��:�s�T���3E���[��%m���M���i��{^�KM�yIC����|?�Bɉ�Y�d)�b��].qt�'�m.�[_��'0/�!a�2X�c'1����w/���ё̟�`���wl(���A��^����薕�^�2���(��B=�P7��c�s���ZP���?l���ƾ/e��iU��2Lj��,���]pD�F���ԊM���` kY�g��5��'~ܸAx�5���jG�ڀ�*�3�VzD�{�a�ʜ>��7%S�J�F�S����o�Xv����K�IHA����#q��wb� �v�6j��9<�(�c�����!�+�R�˯�xwL�j�"�Vu=U�Zi�/�\��^��XQ�R5�nf�=�3��_��7��ܲi�ukg��}и�s5g	��h����?ɮЏ<�O�Ľ�^ %�R��.(����\�`.�0Ր/d��5Z
."��ۻ�tmd0�Ll�MJ��t�:�+Z|X&����.#��P۲�b7"Q �?��:�B�cv��Ja7���T;r��m� N�'OV�$ı��F\�>,SF��T��!���ۺJ�a��S�@�ʔY?����ۂ��N4R�I݆��[�x]�M8?LN�'�߰����^25>��(>;�����쇏�wzZ2" ɩ�ʲƗ��^�)��#��3��۾2�Ɛq(�IW?9	H�!��xÁr�-�O�b0��oL
G"�rX�o{F禵��B�6�b��ve�`�0i�<�_�!.A�?o���xJ)�H���SكPg��>8�ƶ���ɿ:� +^U����ɬ�\�F��9��2D�g�������,)j� T{��|~��,��R�ff���Zq�X��ȇ���;�$�W�T�z�b?®3��.-~�V%�R�5A�Z<��u�?�[��԰H93r���g�/(���P�0�e���@k��I��	���VN�[���X���IqY9,T��+W�|���P�BM��`%.��Hl���8><W»R�7�k�6q�r&5���n.�M���?ҩ�w�Z�|��[fz]�ֲ^����(Pː���e60��`@�u�U/��'гR'b�\���C-���oDU0~��(QZ6$�#������7���]�Pkt�g��o��`0t�a5}�V���dU���Y�s������8��r	]ѥڒ�1~�*�����a�yiw����	)�u��,��[!"��^,1�t�\W(�-RM�Ҽo.Ƃ�l>p^�\��ؙ��
R��<�!���D�������*1(!��7����,�b:w��b|� ^O̼ٶ��)6)��y���lG�)�b_���sv�	�n�g��cʥS6Ĳxf
�qO�o
`�֖r���t�ۆP��)Gˇ#��ٗn��.( Ȕ��9�_B�G6{����`����u�*���n����/�Qy+P���AVfg[2��-s�K1���9^\�ڮ<�����ѫ,�P P���>1
�fB������{��ݢ��@��;�!O k�v}�Ģ_aI\w�ɯ�� �y��GCҔ���s��r�@�=�\}��y���g�w�ͻ�m8^&[k˵��+�~��k2��3ͻ�=�y&ϞpYVv��&ό�i>�#���� ���C���Nb��w^�����}�k�xl�Q��E[���<�<�@JC��5�#5�Gə��pwYއ]|J��L��eڸ<ӑ�nE�ꐫ����g7�ht�=���g��h��߶��b��pJ�fH[}!��1b���4O��DՋ8L�J�6[N+���*��嘮?hPn�BxF�$�ĸT���AL��u��Ե�x�(���S���NI�,����a��1�5?al��T6����=wp�zIDi֥�����MHd��W����A}a`k��f�}���w�"}my�G�r^ݑ�ƪ���N�V�0v5n`0Ť��k�Y�h���/��ut��.�~7ӌ�j�6�����J*��U����!X�6�="��d�Ȝ��`�]������3�Ȣº3�g$�}L���Bo��}�e8r����|2�V
���H�{�x�#X�7�����C���K��3{�;� D����j��C۔-F�N��1fg�b���P�V^������H��t��� %K����t��<�ZLeG��C�:�Fx�%q��=ip{�8�{�P������^��d�q^*�G�+z&sI��W����▷^ ����n�!gb\%FY�U���!�C��������A������\���Yk����^��!	>�X7y����>�XrO ��S��9\���>g�i*�{�i����3SMq��u��]�V$hE��5�Q�Ϊj~�5�2�Gb\��O����V�D&8�^؞N�!=��$�ߊ⧬�W�Vd�ܭe�W���ۚ�40R�E�(��:�˚6;�(j-�(�|�������m���If�T�GF��2���y;ߐګ���S�hJ���0%�=����@�����twl�pX�I�+h"���(�ߥ|m���A��>�q�j~�/���u��%�`�u͹q���9�A m�(s��ux]��Df@T���&�	O�����P�:q�ʂ�N��}uu��+���~�8ж�B֌�{ym��@|k��p?	�n+hD����=9W����̌�2/��߾�s���������[� �3
NJ�P�:L>�>� (6�=4����ƕ�Fa��ܮ�D��$�T���H�,��0
T�?�����U��c�<��7�ml�Xy+9Ѻ��1��`��m�qќ��Aj�BIԇ�rh�)S7oW��i}�싑E8L<7��
q���aF �Uʕv���F��l�Gw�����֫��
����
b���8�խ�E���� y�6��r�l�]�6�JC�[�yD�v�2�<�!})΂�>�$Hȿ����ëTK�� }��פ	�9�-��|��2�Ps��x����m�7h�R�)�����P\t�Q�!b�8��_�3�C]�'��D^i�}bA�D�j�tH������"@w3;�Ϗ��u�|Gx[�Q��@�uQc�X�I#zٽY�����j\v����B9�@�/#3�JD,�)���B6b(��k�P���L�ҙx %�*2���6*�2h"ӰQS����C��)�#��7}#3s�ǞkJ�]��E٬�\L�9���sd&GC�� �;�M��"&\}����Y6Ms�=߯z���/嬕����������f �����س�S0�s��\�>��'��v� ��?��l���+��~��t���N�����2E��Z��\�k�=�`��/��'��)�/�v1#ĕ�;L���F�g��<����u�>'��'��?�l�k��*��~��bEa9�ϴ|�7�xb�\�-�HOh�����r�I�(����9Q�i�!�A�Ԗ*�K͛|�nn��t����-G����j�4ǧօ59V4��%B9��tT����x�\`Eʿ(��.�?/�:%�lĎ����GJ��vnn|8ʮ�}�]��M��ۯz�¤�k������'����Nki`^���w�Q������B�JE;[���D0Iο.��g�m�y�~%z�����U�z*{�F$�*��~�)�����&�Y����Vd�sh����b��售U�2,8���Ϡ%��g�g]>�'�(����x=w_����֒�`�L���V�����X��9��_{��:S�f���P�4�U}��0�(;�*.��~�sZ;��Ī�ο�u�i�8�՘��,GVT��eE�����o�Q��o��!ehb̪�8
�ڒx�n��r��G�h����v�q�q��ϩ��: "�ʓ�����X�j��Z�*Q�
��0	�����2o�WG��1Pݝn�n�Չ�!������4���\3�k���YJ8h��*�������1�^�3
+��s��r�W����_K�����ı��i�+�?z+�(c��D�5 �*��(0��������7W���q׸�h�;n_���k��i�+<]&DN�ֻ�|�͏�]׾�)'��Þ�G��K��6��LPĝ�wQGD�x�k6�$������#
�(�Xu�T��G�?o���� �����2����_�i�<�&�����,�����RK�#r��X����ґ���S�uEɱ$��Ք����C&�>
�L^�V�J�ek�8iз����\|��N͕kݜ{EM����RKd����PN�Gt��V�����g୻>,1=]p����o�㌺��k��7s��瀛�����j�?PK   ��X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   ��X�w3.  )  /   images/b3ba8064-1e10-4daf-8b84-7882f41f3c09.png)��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[pU�y���s�IWo	��� �S�؞���#��y�8�L3N�4ɸM�N��#�8��8i�gܦq�&�qcL1�����0`H ����+�{u_�����+!�d�+<�t���Ϟ��������=V��6)̲X»$�T�+d �Kp�7ճ��t1����#��
9j�g�R�Ij�ӏz�G�Wh�+D�~�F��
�
�T�sAz/��v�f�����o�:�ƅ��\�h���aj�[�>���OSE�i\�A�6��utr��03^b�Ŧ��QLbm��n���kp0��5e�蘁�7����uuĸ�ֹ�!����9XR�1j�P��[͠��ZZ�itIp��=>�I�X!����T����=��`B�����&>Q���!S�ϚR��n�VK��1��=9`j%�����WV(C\$T�_�iD�}� S�9Ȯ�Jm� J9�1s���e�Ң�@ذ5��\�ˤ� A� M@P=l�Z�M�B�d^B�$��%H�4m@x1�P
&��/�F�N�	C��+�H�Y���f��I��BQ?D�x���$ݧ���iǙF�
y��蚗ka�J.��%�Gw��8�ؖGL^��n��χ۶[���O<�ܪ� x���(A�{��T`�=$U�x��T��a4Q= #0L�Y�x�f�A�1,UGZY����a6��a���ӶhƉhL2	>�H�$�X,���QMk O�4��Yԧ�c�TO�3�D��!mx3|�i;aZ5D#�,��f8J5P�Kwbn�+qO{	P`OG�5�w����k/�M�X�n>�կ����Qly����|����ӂ��Ѱ�&mӮ��Y-�ȨE�K1`����#o$R�t�$T���5s�Շ0� ��%HZ���qN^G�u菜C)ڋ#�Z ���V�Q�1f� ��Z��J�	6��\��Y��?��r�ӀaR���g9:�@�2��_�Ŵ�l����A�$̎� ����@8p��C��I�mǍ��:�̡�H,k��"��HH�M5؟��|(�V�R�vǞ��m{��W��L��q�8d7���q~|\xZ��D'T����V��ڠ�(N���$s�8Vnc�$���럔c<%^�u���)����h�,����������-�Oi�Xяg��NK�s��k��M�b��Z�&l���q�{]�M�����~$h���+U��x-D�\��m;\��L��mUM��Y�\�qhh�Q<���ю�Bቲ��eq���H��	M�$���<�F44�I4.]��$���������eGkN�Av}��7��Ň�~��@��c+�QmXlE)T ��!�΢7NGz
����cvhL�3Ez���m�v��፷��~n��c�*u�^�� gއ
�4ç.B�bv�E�._�N\Fu��
��\4� H(�������0��^w��$,\z�M
5�B��j��a)���#�{������g�{&Z�_!3=.[f��)�;���M�����P���6o��'"��ԗ$F�hy��:���]���/�z���sd�#�c0'�
��L,&�� !���@�k^Y�7��֊ h.��x>9�����<�XCćт����i�g4��uQ\`Ǟ�"���v���nBUm-�B�M9wQͳ�_n�P(��X��Ξ;�~��m�.�8?%��$�:���W�S}eT$3k�3�S?�x�ۮT Z�h59���  qCt!�HQ����7$���/n�!��qn8���ӄ3�c����=} a�x�����*R�U�$��d>^�O�:f�bCr���l�����XՋڼU��'6�4{��u	�7)���2z��oW	���%BX>z}��z�7�ϭ���w��-d�y<GY&P?�#gn�&��x�@͎3�"�Q��ߧM�Tf�&3�2g��^s�j�t��m����Z���H&�\��&�H`dd�`PӤ��Y�q� �W�1���pGk�5d\��A����a��l>ч�Q�g�6-��iž^Ы��L���[������s��e+5�a�(k���D��!�|S���?儑&�&*���H8�����۷k֬ѫ��p�Bl߾���X�lR���89K;�؅"�va��H1�|�
n�հ��=�w��k�{��vꇺR��A(�6?��[�jn��d�z �k�/��Í-ᙍ���x�ҫ	��}��;ެ�͋g�-Z�WIkk+������bΜ9X�r%�,Y��u�]wQn����p#��vqi�K��lF)\�	I^!y�S7��mX���o`�|A�<���x��A����a���x<a&3��;؉ža�M.�BY���؊N-=|9{�"�?x��W�k�.�z�ڄmذA��ѣ�����U�p��y}����p�tAaqv)��\�$?���5͓�'Ad�����Z��Y��I�7}���Vy�V�$�U*�l�S��M���Fg���x�5�(����Z4�ch5��SUX�h�e��%�k����?66��Q*��s�N�b���144�MW?.\����a�CFGG�T\}��>�eq���h|�N�ܴ���xЇ�m��&�X8=��um	��zEƚu��|E�]�H�u)�|�b��#M?�$��Ժi	r����x6�M�\g�%x��k�2�s�� 3���~`` �PH���i�����Ŧ��,ߍ[��a�#���΢����:ȇX�7X |1��K��B�L�IfU�^]V�J����ɵV��N�M��gSk�w��^9�a'=�|�X�B3��ٳhjj���l�[�Z����_!cca�B�*iRCR�O�7K����)dI86)C��Q�!�Oa�f>jcuؽ�9~�k���01h�u�����{k3a�����F�u�J��ˍ�`��ԷZ�=FB��x�}����.�����j�N�=�tq;I����t7������f�\oI��E� ʉO��ʕ�+y��(!�{�x�������PV�
������|�x���١,f�S���I��^�L����������[k�� ��dƏ��÷�dqa�5,���qV����g�� \��X���a���D'Դ����\wqo�>��l�I{:��%�埅P���.�:Y,[��<���7%M� j�����MD�*P=]�x%�A�VG(3�Uw܁�:�R��n�k���b����a��=�IN��1
����iFZo,��¨ac��ÞR�F��R��,N�i!��(�q?��	�9=�;�6�7�GC4�"	d��4F����M����f���.�c����J���:a����wMKX�5s��?��yUrY�b�8d�z!˩�$�!�\^';�9�u;�-j���f(<RV|N�L�^�]�	�5���#���� �w�R�'�*@Y���5���p��0�������e��&��Y.�͑�(E�:��������GQ��{:��$�h�ƹ�D�!Q�۲��Ѫ*�c8u� o�����_�ʞa`x1��f���:���\���\Vdƹ,���d�F f
/��h������E���mP�C�Y�8P�ͯr�zC���i����Z!���40�����>���R�oA��;Q�2SO����7:h�m.���x�p-�Ӡ,��`g�ˢ�:]zno��(�ˀ��	�Ȓ�sA>����q�NS5u�w��ށ�ɠÓ�$a�Nb�*Tuqs�����&7\5=R��\����0�̗u�
Q�`�uܩ�q.Kȷ��Lg�ު8:�8�C�pL[����M��	�/b�ʃ�Խe
{Kt�t�6�Ǳ��]��ea��8�m�r�^E��<�hvB ��8q����Ny��!o�PH� ����iE�_�J`�/��߃�'	d�l�ǻ�B:���]}�!�Y�9�9r���b����C:��&�Py�f[��f��rq�4~C�����5���1�\�;�0�:%z��t5�
������1�:�l1�&D���@��ýi�������L<�@0�]*yy,��G�WC�(������X-��9E���^a�t���]j�m�9����,i���;k[MHg~�OB5,��7७[��
�B2�o�@��S�P�L�2i�0������p�|HAy۹�_
g{��Ÿ���/ۻ-eb[_V��磣��P�}�e2#U�����,��?����� �k�y���oߟ���Õ�,6Y�)0����x+�g�?"��,�qqy���Cs�
ޑg���@�NazNS�\�H��KF��-Ӳ&�ej�������x-�L{�0�[>�b�ie���
S�'�?�Pz/D���Z*nmdu�̠7�:Za���#XAÒ���yf��K���,Р���=�gz�$��S	��*
QГ,P|��*�'�FN���9��ȢF��{9����FOnH��W>ԫ*����h���
��F�j���ZzG�z���Em��4�!��4�]sE�5D%�1z'��q�F��8ˑ#�Л��T�4�O�X����\[��b�u�ҥ��ə������Q\�
��W�~��'y��eW靲J>�K�X�;Ļp����a�gހ6Ta��=��>|޼	b�� ���G�e�%�|�݇?1Vb�h�u/�|�hy�ߓ{QO��1އ���Qw�˱B��W�4N�A|ڸ#��1w/�>�-ح:�|�R?����Q͟��UE|��-�K�Z��AuO������[�eA+.�d�D�(I�`s<���e�ڟ���*��������~�����l����~�};���1������+3�'
ٳ��Z�j�:��*�A�݁P3o�P�v�l;����10��G+�N�,� {��lP��iō\K�a��3e�7C�VzW��ho��#S)��䯁�Q��t��63�@���MR{+̆�1�d6�(�pM���d!b�g�������9̭���s�t"1��2���1d�΄vA����F��a�jꚚ���b�R?�E�*Y�-��7v��v��>,��W�)l/���%��P��I�е>+�	�b�!aI��߉���6���A����;��N�[DkS_��������+���'��lwQ����������}@��3~�[�.BYF�{��y�ǲ|>���F���vr���,b
/�w:o���2\犄�$����N��i#��Ϙ����ky�<�v��ौ���$�ARb�|-W�V�p�@?ѝ.d���D��	r�~*��DG�����j�����!��)C�X*����΂wV��\p\�9;�KT�LJ�X�sd��%	clݗ ^�.��я<^��t�p�هwm*���7����m _���!�D������,*?��?�=�m����O������y���e&3���x�b?;G	=�z�p۶�w��_$�~y�|_����Í_��aN��o�6ɩ��s�w�?wX� {��p��B8�����Bj�f��b    IEND�B`�PK   ��X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ��XKm���[ � /   images/e677f489-379d-40e3-bb59-6fe87b8e7dd0.pngt|<�����P�dF��22RV�!BF�13J�>�|d��RV��q�d%Y���>d����>�^���~y�����������j�����0�򮒼&FQ���"�	�~7|:�"{W��|NY���vT�w��X����hk�o�w����������B����۸�?t��wp~�
'��]�ݕ����z	�`8��6�����G�.~�w����A�+���n\i*�SubJi��m)^�.�aaߘfq���M��7fŜo�ç���%����i��^	�H�*Z�2W�����ٓ�2�F}&|�.TT
ؕ� ����}�V{�Jf``��.�-C�)��Yń��1�����t��p��{9���Ө�'�����i���mƱaS��!_V�6�m���mk�_�g��u�����}�f0ms��ߥ2$k��Ա��飵�f
��ved�ʟ2���ffggo�7����^4S���ԥke���G������K(�7I���ٗH��_��'Y��O���s��=0��؏������Tc�4�����1��^v)fԀ��_����7J�����o㧋�Q�!ݸ+�Jf
���g%�~�_��p���Q�^�v���?�nx֜B�G�.� k;���}}@؋��Xjj��N��)�d�Ї�F.ܾ��,�7Qf.������ߛ��\l�rp��l��s��{����,U�7����Z��[[��n���S�U��Ov#�ٚ;Ma9�=�Z�S=44�p��n�)��������c��m%&�a|���rӑ���˗/�W99k�e:�<��W!�~�+%*�W�>��
����j�d�n�ܰ������+�Jx	���z���-9+�Un*e�}[y[�����]�/,,�*��]�]��; ���v����>�sߖ�r����ɓ�Y�Ќ�������CvvV�޿�w���;l������V��M����p�C�ԏ��0������5��o*���l��u���Si��D�����8Qy�-w_z\ӱsvݟ�}���n�g��Rn�җq����zC��W�%27���888�9sF@łL&4W'�񙞏�����{�%�E�ː�'ࢡ��335��K p$�*�ZM����7��~�����7��g_�@w>�쏭��P}6�s��d;�6�,p�.�:�d����^w�L"�	X��sa���Ƽ�˯{ǻ�̍^̯��gbb
��L����g�7�������z�p���ޫ�v,bǔ.��wZ\to�[>���JW���������=zd��``d�j�"Tq��ζ�$%%�� �r�߿o\Z��<YZz�%�x�?*)�-U=��� ��oW�ڎ�1ǋng`�\̀��仜����|�W"MO)Y4�?��Hd��n�t� 	A.T�ۆ���G��3�

K����&IAfk
���|r�\ꥁ�Z�6�������q�`���A���po�&N��Id=�w�v_WEE���4q�� �����T�Y���@�9.;���'I�#N����Ce���R�v�
S�~�G�1@��KMY �~�2<�&y��eִ@��v֊�qgZ���oc@�4
t�G���z�G+ڃ�4���S��D�;;;�7/����>7�����T;�&hoʛ����/�栉S@�=��Z-:�.0C�a��h6Q�ϥ��N�RzAA����L�l����	��[ G�oV��yS�j	F���CQ��}&�p�Eg)#�����#7l���#+���/�u%"N\M�뽔�U�CuY�x�iijp�L�տ��?|xv��2�2f@^��}�}t999��t�Z�4�_8��d����������?��}>���5e��ۘ uf �	JK�#HK�*g�x� ��Hs��z����GW���K��1��{�����VҚ��&����C�m	HJ�u{k��Ͼ��b;�{�$����w�V�e%%砽yr�o��}�\}����ߧ�HhKy�:j�%6'��� Y�21����R��l�w�ׯ_G�TA��C߀�L�2%{`�����`aJ�Ɔk5��m.��6����Ǔ���C���Z��8�i���nc��l===%8	Xf"E�M��͛���@���(a0���w1TDp�z��O���^�:�V^�{gg��@���8xs׏^��U���km-kk�r�d��|���Y����^�s-�PD^�50ϡ�C��i�<%--&�ث�	�g�����^k��]�-�|m�B~Q�C��V��� m%8l�;��s��˛ž�͹�e8ؐJ�@g�p�gkUQ��>�A��	��%E755A h4`hlm�-b7Lgnn�f��Z 4 a,�C"���FӜΈ+=�q�C�{������кdz��Q��|@Y-Ժ�'Gs1D���@[����F����h�@'r��[%`�h X�r�iJ����h�[@$W�q���Z����b�6�x~" ����P�e�®~w9��Y����5?Yi��@��P�R2��Z)HQ�rѭ��{��
�$������3� �����~����Ui�'g����Y��pQd���--�S="�}�2$�Z��y �t�Hu�J)���P����I_�z��6Ov�I���~�&�V�'ˇI��RR���vʮ��{�0�Q+r���]D�~�)+++�R_��1�5Aӗ/�\0UPn�C y}v�Lb�x<[��T:��{o����� ~ ����x��\]�+��ZG�W��$��/��SSknll�Y'�}��T�Ї���e�z�9�p�����?-�����P��\�[�p��p��O^C�3�(*K��������꽵���q�W"viiiOS)`�@�s��E�s�+�!U�d� ��׮]s��Ƌ�-hG�Ǝ��G�|A�w��ճ�r�҂ܢ"��;E6$�����,P1<�:p�f��r���Pȏ�ul�c	��p��s�|�+���p�e؜*�dh�J����o@�
�w��w���^ж�p�xћ7{V�n�'5uuݷ�P��{��nl���^\RR�?[��7K� �UV8�~!=�=����$�X�r�'��/g�+�����Q��e�f��a��r� ���S��9���Mren���*Z�A؂�#�/��������^�X/2؜@@zb�k?���J�JN��0�>������L�q��Q�;�zHt��U+r\�J=<E/�~X\\���ᐸqi� ���!�<����@Bv��|,�� �*���VX=VQQ�����I	���-���U�v������^��C��%�Ѐj;_s�ޒ}���{��'�n� 9H�4������%|���,�`|kk��Hު��]$��ckkk,���hL;Ѐ�- � ]ʡ4�藻O�H����l6\gt}��5m���N�J����!�{n�h8:��̔�5�PS���\�?| ��ejj4���˗�H>읷���\�m��vs��������fTAA�L�	��ö�6Aaaz�fff,n���Ŧ��T6���pv4�ʤ#ww�S�o�h�� �*�f�U �9 6?�h�$�HI� ���悘������i�����%��������n&f�C�d������lPwi�V.����E��E��`c�n������?v�w�����#H;�ΰ\� ��e�n���Z�"�1���M�!e�EB�s�B�v����ɇ�D0�L୘�+ ����44��xi��8&~T�]���k�N?�����F_�U��,��r~�G�!?�vN�`]'G�ATB���7px��HA~�z�	�^�&���Ps���!��2���}�@Ǭ=Yfdf����O�?����x�<�nj� �<���#�����f�fz���i�İ�T�B^��zj�*|����3��ِ�}��_�9��J#/o�� �v��9bbb �J���NN�PU8;� 0�ٲ��0S�=��Y�]��f����7����R���(�V�|bT�� &�i�͂�n��QO��.KAt�/,/GONNB��>Z�j�w��`�0! �ȂȄ�j�D�{��P�}�]�]L3��k1#�yb;vXL�XG�4���ZV0��B������ș���@�r��AF6��@�8s�`n͖�78 �3t҅����O\��==�~�������K��A�cE��h���6_��t8o����f���S����#���M�Uэ>�&%%}xR-]
��₞~�� �C�ׯJt�!4!et"+++!|x��%`&4G����. �c~��^~-�YrEGc�b!|��Y999@C�Ad��A��� gz�t���M����9y�Z��y̠;��J�q���K�佨�*���36�7{�8�9T_�-X�3�" �0e��} v$�'�_��&�3MOO���`��(��������J���Z�Ae�IbQ�k��st£�vJ�+�ea��l�fVj��fx��ƨ�P���l����UG ?!]��� �������2����$?���,�-(L3 ~A�.5�Ta0Ӏ�7� �1��t0i�L�8���	CH���/H���L�ޑ&�XAPR�AK	�YZE&��e����嘸Zͽ`����O]�'do���'�t���!j2���݇��aÁ�� ��в���=��GFX:%֣����^|�}���H��@˹NO*=600*؃?K,Ü���+����f2ek��h�)y��nCgﻀ� O_�����5n���8C��d�/)��M5���0α�~��l~|�����C�|4:���	{�Ook4�t��{G0�)]�CÌ�c�~kl��*�b9��^ו0B�~,p:�����?\��K�Fͽ�Z*�wָ��-��J%�"�xR倱��d: h����G�pe@�C�&��~�=�x����K��������1d0� ������:��u��X�����W7jD[�燶	�{�\6��8�������d����\w��h A���+ >���#t�$�]��_aF��&vo�0�R���-wq2� �<�QQ�hm��E�Jè��f0�����RRm@�A�����$���A+))��ח��
'��m{{>�����p���.T������g�`��9п��ŤW�>���R��8�
�.�B	����ġ�h �X_y&�0�����`l(�גޟ�ɗ�\:��&���,���;�����Z>{&��\�Ĕo'������f��n���Y����)�E�&`���rss� 	4($,�?��&��AS�����z�T�}�
3�^'��%G��_`p<�Z���g	
�\��A�,pQ����Ds�2
b��7)�Ϸy�1 �(g��nm��γι�F׹gsr�{�!§�lW����p��[�'�u�K�8�U�@�y�����#�̠� ��"��O���	��z�~=$Ų���.���`��N>���@֊��}���$ʗ�ѝ�ǅ��ݏ�.���H6�������&�@v�G���6���P>� $>R��+���$��.����k#�y�O�k��g���1f��߄=7&~����T��&>{��Z����ʁ�2m_!�T+�m�[k; � �Z�� 9W�\�Y����c'o[Gn���],[o ��O��\G���1|�c��7Qyf/���7`8T�K��H|��JC|����Sl�!�k�-Z-w�͠�@}n�1�`zkj\�V;��⢫�[��>��.=ƱrLW%����Ҩ�g���F>+����B۷E�TwLP6���������{���dX��QJV`> �͠('�L���=n� {�D�����,j<����`~��i|We%V�0���ĭT�Z���P:k^*!����m������R�������,'_ϥ����J������9���D�9Ch�e�d�:: ��d��5��<�D��!��j�������WK����֙d��"�pT��ᗉ���e<s�;
�-H�A ^��eŦ�w���hw����/�Z�*Ltt��p� +���t��{JP�7 �4�ϟ�j���2�W�`��z�a��w N��{x�Deh���Z����O�"b��]-!�?Wߎ6��7@��R��v&#z��������� g����E�����/�t8g�U6���CXo+��.�T"w�9����/�$��P�q�1���"XRt	6��j����;{U��a�ɖ�{��D
��&��%:M��=�#��M�9~_}�����lɶC�S�!P]���E�� ��L����X!iG���R-Y`P����&|c�Q��İ ��u���u2���!+��m�/�@�������sy��!RPB���Q���K����J����o#��9&�r3_l�vۊS���[��ց7��]fZ�` C���Mf�C;ހ���E�v�`V�����P��ZF~#!߽��
�kr��i��H�Z#(B�����,Rz=����0W��<���H��U�cP�X�kJ?�SE��j�ˣ7X������z�nVx;<^�vH�Wx�d(�s��f ���,�l=:�V��:��߉�艫7���@g��QԮ-(�7ݢޭ�P��𪤞�z@�s�~�b�O���M(�2��0��P-��`c�&��q��e*�災��-���_aa5�Ȧ6����}C�����}�}�H������1�";�b�*��,e��c%K�Ț���.�o�!�<k�5aȄ qx��w��񝳐z�v?��U-�-�#�#��/,u�	t�}9���ٲ�.��uӞ5��'j�.��:�Hn򣋊��|����8����1�Ac8M�Ώ[G�ʪ�ݠ1Pl��=�0��8�D7:�7���1�xs����<\v ��m	��4�U�(j�q\7H��Tr�7���֭��x�� ��.3���q���@9W�F��dȾ���W�$OE�M�R��s���>Ǘ�kl���{�� ��v;-[��Ԙ^@��I�1Nw�U�\Y{�#2����z�$�{~YV�v�C۶K��v�� �6���I�Ns]�6%=���7�)\�����v�(���~����zu��P��'��@�� 
��V�0D�n25q�r�>�0���b�I�4� B'�sn	��������0�e�b��Ƅ���a��Rá#� 7�ٴ�A	[/�5���v2#����	���[^��s�k��)E��e��wt� @�kܼ\Q���6��^���4!:X�ز�^�����4 �CA%�j
�ց�z�Wen�b���XXe`_�NMl��a'����P�W�J��HY ���x��g ���KJ�& <���'�1Ju�����ϳ ��F�=��v����eu�}}}%�]m3ΐ%B_7#7]x �ƭ�)��Ɩ�2����W�����#�3_�J^�Qt(h�"|� �ϚPS�f�Ds~�D�� �TQj��轹t��m޸@94�R瘿��JAû�[���cӈ���@�H�� }�o�pq�4h��������˪p"���'�W�G7����F��աd�j �WHf-�~��V���S�kY�8��p�]�L�f��Ih�w�%��}E�-�"0�t��m����^���t��K�F��*����.㷱��QT܀��g���D	tijB��`U�c�ѭ5�Ni�A�5X���^ph�A>�s���Ň�b�@ޅ��q���&uw��~%5A�P 6�9	��.���FI2�.�L���g67�:��SVY%'߹r�ޠǨ�ac�f6x5�8S���^gL#�̎� Px���求�	�5��	Ze�%�>�l�%{��f%�[�$"́��̐�h���+:�m8O���O�6f�^L+����cHqk����o3M)�*�e��mP����s�ք���f~���MB~�����!�t0������k�U��:��~�w��S4(�|e�9�����G!�����6��l]L���y*f�+��!�{��������x���tñ��̾f-r����E}����Iw"v�����Ҙq�������=h�����'�@>�
�>��V�<_,�
?��)�Z�QEn��:�P�Ї)gkґی�H`���X��y�L�C��)ST����1o:�TQ�j�V�H[�q#mG��Ϙ�� 1A�Q+�>��oA�Ē���&U�O�d�^�|h���(���kM��E�6���sW�Q,./�aZ7`�e�����4�d��L���Ґ!�_��.mLw�]�T�|��;������7�Sm�&��t����~�Ո��@�.�z�ih��~�l)׊�U����rA���;�`����Î��;S�jF�	ﺡ��Bd��b����Zk5�LZ.�p�x�0�ӓu����2�z���n��G+�S��˝�tív#~Ўr�'E�.�89'�,�*���e�@�ʃ�zǙ��1f��@���Z���}�r����ڝ���2��j�\�o
�'Īw!s+����cz���`���ɘU���2�zQ��G��r1��)��Ke9�A�k�2�������J�V;�F������Q����(���fM���.H���3WOj�'�]/�V�Ҫf�����f�7h�=1�٥G�������6�������X���q�f�Xk�e ���bʛ�^�h�(��f}��ȋ��"ۤ�L9�(��� ���ɇ�@���r����i�BE���
�5h�?2����k¹�w@-�,�j�+�^/���N���
u��p�DZ���D}�a��%M�{�j�0Rs��HU���������Zr݅����ӱ�۱�cO<g���A.[��jĝo�z��N�fP�j�oQ�nH����ɢբT�dT�Dro�TS�0�l{�*g�2CY#�{�*&�f�
&�n��>�-0!��D��.h	���L4v1��&�m���x�e�iOB�M���v?���/	5O-nL�
u���2^����t^ut]\|F�l.D1��Bg%_g���z�����l�I���P-9R���M&{w�?<�[SS#(:�*xt]J�����X4v�M��}�M�ۘ��>��̊t�����)��$�IT�Bk6�#@W�t�R�p���X��_΄�1��8,�P�)��Ȳ_��ŝ�U�ۿ�vU�� ��3�iX�y��s�K�$ m��O��~K͛!���7H�5�3�}s3�nU�:7~�?�"�B]�� T���mbX�4}d�`������|�v�
ؠz1Ѐ���W0E�M�d+��{��R�zߞw�����7�:%�ޏ�J��
�^��/R41�J���i�w��y0�#h�h*����jNR*=2W���+�vB��$*�	�n��m�{�E�ᕨ����H���B����Ё�QG> qٓm^V����|J��o⛳>��J�-�U@��af� ���V�-=ɖ��2⁊����0a����UH�)h�&����-R6ɲ�g��-X�6t���G��hd��(�'�{����:B�H���w}�y�d�|)��:�o&;��^��|��U�Z���)�3�'NR���&�_��V,7/B�xNi�aߩ�>���<W+�U�Șߢ)p@��ͅ�q}�z���IFu!��o5m���>�5�����=����Hi#Vn��.���Tgz��U�ҍ�>Y@�̦�KQ��k�ҽ���#Z-��%X���`1G��+T_��O�X?�܄}���n�W�B�}j�E?GI���P���}&��7�:m��_�%#��= �^������?.߿�����>ʎ3p����u0�h�����R�흸,�c=D �ޮ��٢�O������_KK}���ˮQ����՞.ǅZ�TJ$��6��C5���l�H���@5	��L�ͦ��'B�Z*��y��$!Hu�(ްq�da��
�X�.l��\]�~�
��d�X��[n
܊��^���@�����>=�h2;���J��g��0�&��.\�îI����?qBe�?�<� �ɘ�����b��,�����.���׀AeFF�lt��#�D}a���2)�NI �T�,�%�{�"��.�k�
�=
#^�.��W�G{�$~�]/ ���9�d`�n����#q�=���[�pӧf�,/}�����d_�o>~�͊8ć�vyrd��0{���a'�l�E홻��[ҧ���'%��9M�X�U��	�YL��0��/Bt����4��*�79�3&0����s�[�?���D������:���P��
t��'�@���
���AO[u%��A[�= �f�䄡2�[ ��p?��@�Go���`��`y��H���;�O���q��vrr�b�׫�j*!M@���6`27j�>��V��Q� ii6����Pv��,t�s��T�6zv��d̪��~M�����c�%bؤ����UL"�}�hm��7ڕcu��24@��?�C�-�������S�/�^�úΎ475��U�^��C7
&���:��E����(���|�}��~���R�/��u�Su�_���rn�	���$�(�1~.��}���ҧB��n�t����MQ��B��:(�}aU��,�a>~v��[~��~�y�������b��+3U�,�\���J��D��;��NU\9*��	4�#�!e�B+��֊y�x�)�u�P��Ex��/�A�n�tKl��n�pg����L���)>9MG�*����E����+��Gۆ�)�z���P���~e��`@|�=@m؃/C�I�ϫ���mnm�6¸xRZ�BON�?�1CO2X���'���n(�&%cY���{���x8+tUA�g�eA"{�Уv�Ŝ�Rb�f��(((l�A�
ég�X�Ⱥ��� =��g�И�H��#�Kq�fճq@.���L�������6��	�~׽�5��*6H�2=H�gf� u��c_�Wq�BF*9�Z
u��2d�d��_�{"�赫@Wuёl�p���e�f��o������������-^j+���o �>D3�C$׏P����%-$�F:�s���
"��F�A�ݩ��F�Ao+�*H�~0v_��8os��A�-M�f\*�kQ�8ʨ�~�B5���)�`��WV=v��������@+����:0����꩗c�����B�^�AF-�2G6��tτ�ڱm���8��
�Ȳ����
]n�;�
F��"�vu���TJ�@�r��P��g�!0`BOAl�����P%X��9x_?��Z�J����C��2T�6l�g��⢑@_���f�9��u0b��lŘ����	�`@���o��y=((Ⱥ��S	�&'i�h�w�� ����8F�œ` B\�}�`&l��C%:o�h�:�8�����?J��~R�������E:I�*����k�g�H�0[$�fg���̭N6 _AF�|�qv���q�����z-a��y��ۯۏ@8���J,����va�|rA�~�T��r bz���Q�N�P��.���N��͓�o$K���~/
Z�+a�3]����]U�����U� ɂ`}MNN�]����ʛǄl;��\(����_�َ[�żSmp �1"���g��Z����0��2:|ʽ�����G���آ�g�@��(�&	e���|9�繪j?���ve���[��qϋ� ��k{9A�6g�/�랣�cN���[��$]��rRX@Xf�V\AAA��86@e�M��	�R��k���0ϲ%�*��]2"D
�"	��,dA�J���1�>b��r�َA�@��#Y����V���&��mvIj�x%|����W�EY����^2��u���� Zs�^UK�A�@��_B���na���a�-S����6g���Tg���������5]_%a][����&~~~�-[�ܧߺAܼ�<��
P9��V]>���s�0�������Z.z��0�
۔b������2G[��3����t�%�U��7����Ub�+G1�U�����Cb���ϒB�H#����tt���N�u�_�4ܛ#K�~�"��P6@5��B��?8Z�,H�G�?9���P�I]�xI�R�W��/�9�Cj?���R'Z8"�EW.��f���$��K��]x�roa��(�]MǺ�_�|I��}����g��G��_ � jHKSK�	*8�E+;���l��0�7C�1O���b;lLo �����Jl�*f#(�N�� ي|1A���I�;h�5St˭�}b�T����i�s �
��Wf*����\gFe�̊d@0n#�f$(қ�P#T���6���ԭ�z�s+8\��9+)��cX%���C���	��f�����*l�[�:6P:��Q/��*��ά���Jx�AK݅���"�I)��OQ�-���L�O91?6�y��\����Yv�hI�\����X�֡� =g�k��!�����P���i����J��������᥎�Evs,`�����?�\�Z�>���/��X����'' �ݔO�ۙ�^L�Yk�������=��	�6OS�\����}F�w�%�A%o䖤���Ӏ*>��ݡI`��?B�,� �l	��>^QA����elO�]�ʯ�|J����sMSA����A�s���/���M~���OuGĿ�w���Pux�ą��]k����)b�f*1�w��h�#Nލ�ۢ�XL#�E"��r�u��cs}��Ņ�';v��rN��,)vk��s�Fr�3�(�3���!QD[� �����މrB�����R�2�[gihh�Ƣ8��B/����d��\!��t�>KŴ��[�N�`�vp�>�i�ޫ�T�rՍ_�!�7�X��|�#�=�r˽.8ᗮwo��V'�A�Z�sh�i@���ǜO�>u�n�����jFn��A3<2���<5e6�utYF���썛��G�$#�~�V��n��4(�.������59H�Ѱ(���}%��>7�("������ޙ�qN�hk/	�
�K7�����������̌��G#�x����"�I:��_�*�%7!4�O��>sP'*0�Ͽő6��e ?�?�f�����|(��q���<�h`B�I��D(�dĸ�ɓ(��(�i�\�G�H���_�x!Ó����m	���vzC��M�i<b�W���8W�k7�j����n��zqG��k�Rv�J�K�\��Ml��=��l�I�
�����8%���h�{Wiυ�����m!{yHĄ���r����)Y|#1�(�5:��鞐���>4��ŕS��i���c|�l����ߞ���w@b�ӥ~��/"�<�D�vlNk-s�`�,��(ߜ��>?JFC�tt�6ZA�����Ƅ�+�ǡ��~��O����'7�X|NGe��-mB�&$'gefQRR:b�%#���\�T��}sV��?�<���(BWq��&�[��[�ð����<�c�&�>}��z���V�
��l��,� ���!��Ҭ�rh����d%X[666:��ʄ���ZH���!�[X�`d�@�������?ES�B�ԯi?hj/�����W�A5� �1� �r�F!�hL�Z%2Y_x���C@�cӔ��{(+\��i��@?6�	��|@ \e���?�����=8x
�gbҲ��dW�!!$���V��]z=������bs�ܼ<Y}��K��k�)��D�uW�v�n�td�s�YZsl�
�����_&b��Nk/|�̯dHU��.��n#�$���Ӓ'a����İ���	�9��԰��#ݠ8~�zU�ea�GGG�Ci�?�q����O����^�ޖ�Oȧ��3�O�d@�0�����I�J�N���)l������q���^)4�waJ}�0�+Ѽ�;ѱGΠ۠��k�S��T��f���*��^AZ_���>#�bXb�Q�=O2�E>�2+�5
5�)1N~W��׵kr`�����J(�Ql/��q�X�v��իWϫ8��y$H��"I}<>��8U(�;Ɨ�����̕v
����|B�a��k�m�|G����͗�KS�8��{<���?�2(XIF��>��E���3_ ~��(׿oV^�o�5x"�'&/�6�(��+dV��L�������W�M�g�i�C�Z
|���y�OW;��ƶL���o���X�_����v�;����� ϔ���4	���,��D��^�U����g���5i�m�����3Ϫu�B��5U�vX	}~4D�_���[�aK��e�cO��T�������e��yE�z6��)��K�hx�_�s �Q ���%��&y�q�"��Y#\I�	�J\��֟�̺:������k���:�Q��3+��t(�u����r�&:N���r��������_�rV��C�Ӟ�<;�j��ϩ�{�0�3؏ԉBG�%A�@K�_��5�S:���ɾ}����($j�g�,���J�k(�@�1�����ǋ�N�+*��J
�e����z��2S�k�!�=Wa��YaP���  �sL̟�Z9�Nu�"A�K"saU���Ɠ!�C!��o�`�P"d,-��y�nA�m%ꄟ�3dw�*���������Y�Xi~Lt��ؖ8�l��8��/�3D>tq�m�8�t�ۊ.N�bv+���VM�Y��jm�����	FV�xG�ݝ*�y.;;�dD�$�S��DZ�Z*"1~v$���ɱ�ȯN�qg�֘7u�����s��<׮Y�k��WUU���������
m �Wp3Ap��Iȵ�,�od�����|�G١ZU��0��{�][�
��32JĒ�5UU)JY��%��z�1����R��֓E�0ѥz��ee�uu&���H1X*6  ss�?�x��qp����_U�=���YAl�5J�H\�$nש�At�������:@�Qx��#5��%Um,p�j��ȏ_[�ry�5~~--Z�y��݅��ɵ�p�y�x����t�7^v�v�HF�����`P� ����o�:��%#]����VB�샩�͊6��h7F�� �b�%KLL,���7�muuj�Y�$��zz�{(\�j%u�	}��8 ���u��@O�O:�j���0d�u�����OX�YqFA��;K)E�H*����L@U�;�L���ڍ+��I����i4+o՘xĽyt-�7�����EyF�a��!�ڕ�W銵���q� �jc�����d����:���*.�p��:/��9yG@��41&Ϟ��X�u��/u}��o���Y�r���^u^1����x�F�8���%�6Yܨ_���^� ��ر�6�g�n�M�[�f;\��1Di��{*�7�-�DL�>�� ~Bh+�������ʇ��Z��9PV^�`+�f/'�s#:-,FM��5h����M�G,���Z��{�X5� Ԍ=�B;Tdi-�������%׾���7��m
���Rx���xTms�kv����-�qXR��?��S�7~�������) �b(XMf)����<����J�>-�e� �ݲ�6fni�;�zE�E��b"��(77�k�u��"m3f_�����Ȅ<e��0%�?�� � ���ڎO���Su���;�ig.>��GY��L�ك�f��Hm
r1�_��W/\0��T(�Ǧz�ѷ��	Y��e�QR�����İyKL�=G\�i^ϐ�PV�����Ȉ����+J�o'@s��|U�(��W�Ͽ�&�}��$��^L���\4^�x�X,���s��Z��׹�)0�Y3V��ܱ�Ir�K.�� D�o�x�7z�gt�S�Ja�<��Q����.���Yc����!��0��?}������6&{�ѨV����5��0,��谀7�/"o!x��P6���?a�ph���lr���Z>d��8`�JXo�����%��BҺ�UU�tg9?��Á!a�v���޳�1��>C�
O�� ���)���PV�N5�Ӗ\���i��\q�++-u�a��u����5�4�ǈ�S�A�.�!ڒ���P������§P;>=k_����+��#?�����/��pq)d�^�e�n:�N�]� �������/J< m:�zvmx��IHdu-b����A�� P�tu��|,mr�HJJ��'/^m\���V�(���|�,���;{f����i{��'���2��)�D����ֈ���.�y���<z��f��V$ ��ōpm���˥������E;n$��VYooL����r
F����O�Z�	�6�}�㕵A��			���Z�SSUU�����s%��o�\���US*��	q�]4���̇n4q	0j.*J�������[�AK�t�a�QZ؜.�㸜s��òw�J�{lO�N�"��Ă�a9=�sz�!H��y�=����[�>@�>�D����������@5��J�,��=���Z�4����TX��VD-)&��H�Z�[��(�;��C��j�����y����]������������a��tP�'>�#��훁ֱ,���0��QZ��T`q�����Ǒ�/�cw�T��W�$
�^� ��[jY1Y�m�nZ��,�t����9i^��c�;�ml���l�Q�o7��~�V䈐�шy~kY�쩋�#Q�t��!d�r�ɖ�ŀ�Z�'��������1��[gO�zy1GFF~������փ�n�d��B�>:N� ��}�>�ې��s�۲i8G�Յ���������Լ����^�եv.��g0�]��(k���kz?|Hd,��zHM�ﶶ6�_$͝�F�rdY��2;a�����˗D0P��[�&�� !5Z�k �^"�m�M` ���V�������!*���TJ�_�pg�l*L�$3E+ t�>x���.PM����]/j�����{\s캒��v�O�GQo,�cM���������l [&Nnm�~�4{0{�����^Э�(�8\�>����Q\���6��
�����7�= #:��5ى����Mrj��fY�q/{��y�m�35��"`���gc�vsW'��WZfڒ3�������)��⺭�<���56����!�e�JC�x��K.�KN�V5������]�Y�J�U��J'Ѵ��>{�I+JUFF��޻����=U�00��D�oS
��Nۘ��Ά�^f�u��=+�dMo ��������b�ʄ''?,˼͙^�?m\�{�����u�0�O8W������	��������zFF0�0-ON>tuu=�\o_��F���ʒ]<G�V��rO]}�Xl��x�Q̢����㺔?��/o������W>Ps,���2	�\��k��($�3��[��DE5�)���SRRn���^� ��;�:&�
�wY�ӧ����y<�B��C!�����䍋���W^&t��4;D��
�'�(�fd��
��`BKK��7�'��|��<R22|��n�)���"�q�{���[��O�Lk�j�f`���T�-Gܧ�V߼5��k\�_T�S৯�`���`$��|��˞�����}U��n7���K�˃�>*ٚ_��}��2�����FZZZzH�19�����asf�L~��l����ܯ9"RI���]Ns��8��E���x���f�Dv��s,���
����c.n�8,96��5���zy����R�f��^�ab"Pm	����ӄ��%	0�mwx˭垪Ɖ��~��u��,U<�%�]F�~?Wo�Z�ܡO
�*{��~��F�q�1�CZ�a�m���dـq<��
�.���\g�@��XR��!�A�'�ݨ��@��d�Vb|ϯ.�j'/;�D�`��b�d3�������h���]-vg�u0���+���?����n{�A$��F�C�E�iA���C��������f��R�\x��>�}�r�{�9�x���9��f����ϢAX��r�w{��;aW}lgL`�.Ilj��.z՚�2��>�uWp$Fl��Ԥ��d��G�'x:�
���#[#&~ ���$�>|�0�BFF�=;��^������;e�c�3M* �/��.Kf�JFgffn�������Z?F|P�4,��k����~�=[��P`t�൏N�N˹�P�׭����I���>��z\�9�P{[�`�����W�|4�|���Dp�g���DDDn�ME�2
����
(�����:��bl���k���%ib�IH�T��^S �O�5fv8x�A0�t��OÀ�XF������fVD��G9�,,�ńhHi���=h�d4������X�1���fim}�llj�v�}g�2��ގ�W��������X�#���d ��MQ?�7W�39T�
�_��(���W������	�	p=�l��W-wW�d�f��m8r���jͱAAE�:�l{�!77�ֆ����'xXߖ}f~��3�}ݱa��9{�_��ׇ+�ˇ��j_BXW�~#��Jθ�
B�����f4�
�}ɷ�WnJXF��9�܉Ҋ;��=��CK^��H��OB;9�(�hk�nf���Dº2�cZR�Ą�$��"*g��=�J$����jC�l�Msϵg?20nes{�fd��n��d���|ˀ���ᡔJ	�T��S�>�]t�﯐�8����$�ۆ��I�#p��af�oS�q�ё���>��a��m3������҇�M�fy���������u,�9V6tu����>*M��"�5�5{ssx{�/A��C)��ɬ,�z3�ĩ|����+�B;}�]Yvޜ^��a8'���aP6c�{���e\�K1X�O f�<N��4W�����gK��\�݂�
��͎n��u��R��5M@@�=� �����dT1���!A�R ���*bg�><���י�{�I2��r���D�4T��̑ N=<<vM�B2m��9�bc�57�H�����d�@R��o�	Cqu[�������~��z��m�W�`7>��,�:f^�=��q,bT+Y�`rt�uw�S\cs�����j����l*K�V���>@q���X+Y�S���H�- ��s����wrz�$!�:d �7�@:f��a��_�qhih��ˣ3��T��À�� �#��gA�@²�[���\��NA�ۘp6����p}gH�|�ː��O����1�׈^�	^�kkk�w��;C/b/c��n��9�F��a�K1���'a���L���$�������(�,-�k�߈]AkZRR�����EEh ��JKK)��H/?-�����/�=\�@��것]b&���v�� ���1n�����������,O���_[-։�����]H�G�g��:��h�V�����m���ە��; s���u�QDkg���q�,`h_v��,"\~y�iZU%�%k�]Cj������A�v�歹�U@�r��������)ui�\�~`��'
��������9 .��� ��s5\�+]4��o���<��I�/*װ�X7@�N�G����S+Gߪ��
O
��SUSSPT���$^�%!!Q4+,(05;*֬)kn�h��|TC.,,��[k����l5�Ȭ�P��,��d��!~J�VR\,���2۶%DiG�R?6���G���XF�g`d
��}�hF�	�P���ޏ��ZZ_23) �0��=S<?Y��o_�מC�u���p~�|�80 ���Ի���䠟�����Wu�F{��ºR�_�d�Zp-_\!�����������'���_�����g�1<!��jk�e�p:;;mx����������������	��(�E����g����߂ݧ�������C�و����1�R�X����-���d���)]/�!�+�פ�� ��[n�s?��tv��OM�Y���2�{9c�����T��`$����.����v��B;�gg���U4 �n;C���;0�>���`a�C�K�͉1���Yr��v��~D| ����|�i^�C��� 9��U�PxD<d�%P�44P���'u����M�#�G��o�������2o��,��@���������!!��3��&��.�mt��� "u�X?��W�F����k~>e�kT�=Q^C#dtT�V�$u1!6�ըB�3]�j��\�{M�w<�]��>�/g�B�t'(�	�RL"��EE�%�jJo�$(f�a9 ����KiYY}GG��)��T�3^q��D��ټ�r���}�E���b���9�b$LT��0�=���a�0����`������_���/ד�<���7��_��]���'Z��OX ��΄c�d�&)�g��B�����7�����t�@G�jX2�Ut��䧺v���no8h�;ރ��`�B ��<���TWӸw��̡�ML$�p_@A9��\J�ZPP ��J�����fv"F�ȣ���	}U;����z�������Ȩ\ߧdl����w\�����+]a���s��=��"R�OH��X*�Ce`d�"���3��K��!�W�}}N7W�r�H�}��¨�� ���0�[R"�븧�]Hީ�?�ϙ�*?|�� �tC�L��+f Ƶ.� �i�QB4�U3�hA�m�6��x<4���X�~#-����G�3V�k�zN�c��g=�[:��F�Go6_���,.�νeѪ���8qrjai)s����X�����ک��Atr�0+e55���?>��V���X]�>$a�֛gg��؞WZ�022���	����9�,)��6����� N@bb�/KP7�>��vB�]�|'&�r~E`C����Z��[}l�X*H���0eG~���eddx��Ѱ����|@�7��4�ڴI�����nڧ�����u�g٦u�f�岗�<1�5k�6du��';�v1��������''��λ.{GG��8�^��n�G��
M�U�?yBhs���+Ի�I�Im�п*��q�����s��IJ��#a<Atܫ�xh�ϙ]�z]����LtYXБQ�6�g����Z�"J����rh�#y��<���t��,mwk�U�-:�v��VU�D��&p}m[����/_���?����
|i<��N��ں��x���)MfGŌ�(g�9�f�U��gd�7���ZY�bz��888�F��:/.x�����`_��,��V[KKKKK���^u0+0�)�?ޣ������1>�;�ҽ���0��f����e��{�k��G�d��Jy��|��y�W���>������u�mX_7�*�[xi�� k��@M|���?�/b�����8��6��G�]c>CF'D��J@��9��,�s��M�G&����g��䋠�0��fIC��+�:��!���͛�X��c��p��HV5�5�^�	�U��"�f�`�����Z��]��m�}MN���V�'UX�q��vzz�?�U���A�ؘ�j����E����9N���E]c/H���f�p9��2��H���-���)���I+uo%��^԰���7��?�;�z�23/oO�C]II6��E���Y;V�monJJJ���������xl������M
��W��oVO� ��H������J�A,k�n*��r����٩of��[�us}MS=�_��pa�J:�i4�dѶ�6Xsoo�L�X�LNFF��A�f%G��4��0��NBS3�r������=����cK'�@pS�f�+���ѷ\���ŖϯrƩ��UOU͡�P׭�-h�&�V�m�TԼ4WT衒{sMB1+��M��E�x����̌a���H����{Mq��E9�3/���?�yV�Nbբ����㲆WۧTJ����9E-�C�p�[Y�����Ydȫ\K��dw�P?�R�.q����¸��]L^D{��p�L@�Yz|jZ]M
�*�l�E o�'��Q��&�a}������ޜ��[N��Ni��d[���#���}߂PՎp��=?K'�����Y��Q�W�`�X@@�nf����� �h	}�ind7�b���t} � �uq�'�|Z'�8¥ϝh�P6#\900�y���l�����+|�:����J��ۓ�b�ѬZ�Հ��e�����Up3��0��L3�cBĞh���N̺Y��߬���}���0x�:�	��������T2��p���*�O�`a6v�̫Oj��l�ԞR/bz�#q6���l3��U%��3,/��"@�6l���I9V�8ɥC���Ϟ�Y頢��'926F�â���+2;�CDDT���������=R;8:���B#�.X�+55z8���L�j���T*bl����ԩ~�2b�[��������8_�D�jhh(��V���7V�jƴ������2�_�h�!<JG������vU`����A�X�'���(?�c8-;�j����}�IGfD�\Rؿ��\*9������p��&��"{| ����ϟ?a~��S1��xO�;�LLB"8v6q^El��v���QF����ً����s�;�CY�R�7ĥl��AӞ	R���]��̎�h��Ƶ�>H�Q@A���_wǿ=&'Q�l�ۨb�n#�o���FQQ�AY��ڶ��Jw��BN>�P ���v�r�d��'�Ǖ�J
P�	�R3f1��s��Z�&��g/�o����51��^���s`xO�n��
&D��3}tn�;�BYU�4�1����,����~�
�=�s�D�4����!gbp�"�Tpp�/V�,��s&���6䜉f�����9-0��Y��Du��	��7�PGk=��dN�
I�����.N�[Y�Kc[W۫�y+nR����41sG�К���\����L�)-U�J^O���Y]Y�����(Gw�d�}�]ǆ�n`�w�Q�?y�C�s$�9S�̭-S&ff�݋l___�[��U��u�M��LLL��ʨ ��:7[ҳ��sm� �^�7AWo@�5����	��Y���i a|<$�Y1�T�n���a����T��#y/5�����y򚚌q���//V"��(?V;��緁�r�lY��b��
(&��9��#M��! b�.�����n��-kEvҶ��A�\?G�oIikq�H�mIc8�<B�f�%	Z$.�^OT�y�w0�"��W�#�>���ui����N},�˧��S�A�y�X��I�f�@���I�4԰�ks�{�?t8���B���Oj�X^_�ƌn���Q$JKb�ɽ>B���'��8`�Q1$P8'D��L1����J���Xr�%$�AMV��$_x��B�! v��)����Jd�K�e���z����K��Ͽ�*S�����])��}� xz��j��$zg�X�p���v#$�V��Zڞep��m���e�#ET��M� �h��}c�D�}�\ ��{�V���M!y�$-�8Y�oϵ}ǈ(Q�����#��ǱR(��������#��;��������c���'�ˀ�"aH
nzh���:��%�k�V}����3��~��� �qM��f� ������<Qe�GC-��{���B1�O�$Q���޸���Ǚ��ȅYM����1g�?:h:'}�/\�ڲ�j�;����F#,�����q��|*
ߢ�BPK��A�"�&`R��~AZ��	ހ����Q����(�^�xBK�t �&�'
�rZ�����s&Y�"^�y�"����;z�0�PYSc�'��5$pUT��̾6_g�].�}�)qhA��:��j?N
�,E�$������@�+�[��Du\:^:���|?#S,�)��`C3�&O�ǨV�Y
��F��y>^�J�r��]�"��\�f���e����pk��$ln��hrv�\��Ĝ~�gX��@�@�^y�B���F�:���6�ϛ�~.�	���*�{�����y��Vـ���)*)��� ���c�;a��fF�A��؄"U�4�?3��_����)�Hpv�x��GQA������X�����>V�ؖ��zb�ȗ����&�;��	��r#[Ǟf������zh}Y��藑+"�������.��j7r�b�>c�>¥i��D�ܼ�����Z�5Q6�\�����SMY��LQU����p9 �Pk<��[�ͬ��n�&%a�q��l����BBF������᭲N��X�Kȑ�����ίu�1���8�����
pG��˘9��r)<�Ue����auu��B뙚��f�
N��Wl||���A
r��MC}=�R�ס���d-��������@2��O��#�?r�LO-//��p��%LyEI������ї�Q�ի��`���g���G����27�td��9Js��$���n�E@��+��o�l7��Cអ����Ihrx���4t�7�qs{�a��D�ʸⳫ��F#`6b�������n���ut�>j����4��'��W�d�3<ȝ>D�����Nq�Ӥ�t↛7��JI�@AI)&f�z��%0���~��\D����[)��z^��A͚fd�y8�����r���}1ް��\_�-��C����ڍ!�흝���|2S�G9�Z0��/�M�(���a���C=ManT�(Ъ(�78G����d�!7�!��&bX"
��%��=�5m�E?���"y����v=UC\Q�8UYss8��T�#gb �Z���̵�z����C��Xf����v��ڹi������Qa'p��
��,��K{5\ykz~�z�I�'|�p�����	N03|��Z�k�SB| ��}��h ��":��Ry�' ����q�'��]:r���$����Ye>�79@�^Ⱥ}A���N��I���ˬ�G�C��nr&�3���"q�O�ɦ07::9q�b�b���Ց�Qt^	�.��V[W�.)�jh�к�27&��(*&���g,Km�d?�e�c�;tm��Y��ٞ��se�UV�b�����c��x�3M�O;�ŕ�Q���M�����}Z��.��~�vVT�P��˗/k�60�'&��}��ʻ�|���I�UVV��1#^EEE1mL.�u0����Ҭ����h����@�xk����͡����SA;���'G��OE �����<�|��H�9�D0u���b�����������|\�vMH��86x�%Jkv��(�l�6��w�$����ks��ё�f���P�I�K�1H<z��t�Y`@@�%����K2}���niրW�FM_��y�V�Ã_�%!v��הؗ�OAc�{�41=�d�<U%�)Nh�a����x�w���O��۫�;>�Ka
���A>||�V��2C�;$4JF�_^@��D�_�4�¡#L'^(3ĩF�lḄ�v����tP�|D����?��R�~�[VZ�[K%%e��ЧHa��99Ԑ�9;�?c��0�
j�=A��{�B<���	�T�r�_���z���z�$DfA�?��C�tzifVֻn��{^--�M=޶O�m���3dO�iJ�6jT�-((���%�������?�r�����jMޘ�9B��Kw�XH�9�a�`!����k�ߴN�[���8cxq��Z�ǘ�j����$
_���RuyX&ȫXU��K.��KN^I)���оw�*ߓG��e���~d�)����º��=*B�AЄg����=�%�~�ؾ礩��ө��J���$M%�B���6v��������aӁ&��I�Q�	5�[/=|����&���"����{5���V-���z��I_����k.}ջ���@e������ވ���ղQ�� �לA���h54a(���V����tą/������UJ�_U�����@h�\t��qr��)�?215�:��5ZxP$��mמ�b$����P����Pd����-}���k�8ހQ�Db��L 	>~���&���r�%h���@��G��`n/4�`,'U&LO;"��?f+��qFP`/�N銽&}��49$��I2���ŠS3����[ S����+�0��qqq�_H��R�>��x����� ȭ�)`�n���$@�+3��yh��-ų�����WΪ�_�<��V�435�29V^��u��'$80~g8@���,ٛ�JUMA��I��6��|�n��\�H�U`b�+5U�c�L�^KsSӑ�,I�h�ݡ�c�I�KPM|x���?p�c ��>��P� ջc��~75x���n�k����O+���F�0��O�ǧoUUUm�z��N�1�ߖ�
_~/)��>9<d[p?����{���t�}� ���C�0X�v�6M�ח���E]���w��*Niii���nhE�[?�3��5ċmx�vd����_E,��6�C�L��7��w�\b7�� ���ׄ�I(,ܰ��x�Io%��|�^�e|n����g�d��g�^�s'��T��k�쀎� F�o*�g�>3#�-��C�Q�U������/������Q;�@6�u\�>�|ft��(Tw)�v+�����㛗"��**��D�]aDBy�j��`�c#�����g��[���i�GB{|�A�jj����,�]��H��TQ�<ݙ�g�����߿ه{�yyy�&x�@a�G�D���O��x��wًg~I�0�ٴY8�.3�����y?����i�d3N��N�y|��.O�n���h	PNtuw�		����:A��^�5�p�N��"��6<���V�k�A�ronX�/���+pR+++�f��55j�K� f�҃�����m��o�����k�~��v�T�^mm�C�n6��o0������J�����&��U����-CSD=Q��Hu�r��QUU%�tr6g���J�Y[a��X��6�k����	$����^���_���E5�KR�T��#K����m���������������5�'Ph�hk͓����\bnA*����	�hb��@*����{_/Y��55�n`����>3�q���%��Xl.{��v���v>κ����#Z��m"Շdڄ�E!��u�#��qp_!Zl�i����:�q�՛7]%�AZ�;Q���*f,��"�S��M?dֆv����y����Ը3O.b�����+�.̑�9~�JpK����аB��n5���T��"�2+�uE'��(n�R�N6�Y��z}�:^M5�"��Œ'\qE�D����cYn˒T؏�|�7R�Cu���Hr~N�JCC����Կ������ȧ�t�oL �;i+uh��'�^�,�:C_���GXă�ޠh���n�!�/���@����]#�D�	�تR�����Ͱ֒�����""�oJ��P��ڟ~���@ɧl��͒����	���ؔ�w���s����>|����q���3:�q�
�\=�L�M��*�@Ӄ�t���� #[]QM8�5Ā;r��-g^�8��e=�h�3���ɚk�S`���Hʅ6�Q��w�(pQQJ������sͭ��|1!�и�ҭ�����V��0*suw���0�f��r��%����h�E����/ i���[��C�����x���Y�B}�ߦx�G8T�"H�B���̞#]H���c�?ί��M�Yr�i��*���=+�PSS{��EShÓrD���8��TP]��.пf�\���A�Ó(>x$߷ ?���='� %�O��ar�8���	� �ݪ%;;���#���2�Z�����+�J��:G��/�d��T� ����B,s�T��ۍ��""��\�X�W�l�e���% oL�;CÜa�:�
m��P�
����%J_U����E��H�=�Qr&��{��Q�p}b�C�s�U����/��������L�l�K�u�5<2�ag��,��6�>������x��S�[Uk�[aؾ��~�r}NQ�WQQ!�m0z}��khh��=<,;���d1��'��J-�11����@7���۟�$I�����Q��w���j}��C���ē�[ސRq猈ά�H�R��K:���3�0����-��mL&`J� W�3�JLB�g�ttTi���d�ǧ0D߶"�������yi�:S�+��F���Cv�e~����O	����(5����H �ͬ����W���u?lCV|����	�x�':�A��?ZwN�a����݁>��^������cu���XZU�Xp�:0(���O����Ķ
��t����-���@}��mm$�:Ob��a�������]��S�R�]?�;�8�p|0�0�7�B<�Q�dU[n�~�����*3KԻ���x�OC��BK�A"t/���2��`a��S�">�q��K�FKʙl��N����^���s �?��6FH��H��BCC�o/x��`��w�x�����*��;;;���  QGa�����5�"�~�9�������Ҵn�nd��2`o;8�88v�7@����Q��$oV��;��bL�m%>}���._����;�/1`����F��e����s�Qm\V�s�� �@5N��ﱤ�?f�� ��/N�/ޕ%��"y=�ʙ�p0q܎��I�^/�Ź�`g���P�mT��+I�h_���'(T�]�C������.ЃG��e��g-�>3���{|�����()�a� �Bd���{d�L�̠�k@�xd�D�%m��Oh9Z�s�.�
�� )M6�)}FRq�F���|�D"���T�.��V�S���ݝ����&��ށ���QE����z���'�ڼ�077wts�Ev�SC�� BZ��Xr��Ĥ����G��O��̐g��Suc#��"m����ϔ����{��(��4��+������Ν�:�7����$f���67��X���/���Y�� �ֈ� %r���a��	�~7�f2>+���V�?<u��dޕ~�#�i*Z`�bx�"off~1Vz�+C5��M�mC��ą+>�G��1�xި|�$�����M�K���G�G��jU1c��;�pqs���C�)~�Vl��:;��޵�1�e����-j���vX~>}���T	����㽫�;@�L9gz�LL�ot�o�̨CQZ����E�c�(��X�<����z�����nR7鄩;1-��g�t���.�0ڐɄ��ά���O��Dc�>������u=-�Ԁ�z�.�n����g�rh    ��Ud$���_%�Y��!�h���1zcf�������v@)?6r�p��_PӴ��؏,��'��7p?�3�T9�?f}ty�^C����l��������K�0���~_�>�)�ѵ?�z�g���	�#���g�B��2�Z�7�AWx����՟���x`�3ӹ��E�%pɅ���ąD	%��|ɘR	`R�\[��?ڷ�w��0Y_�X�YĘ%��~�%�J���:.(������gf{L^'�h�����	ی���xm�6وPo#ˇ���4�c�hp��_��٭�+D�spPq[)G�e�E0�� �+!�U'*)-�QL�#
�/��l6��f����T���%JҀ��&$$0���yy�X̔�H�y��򨞽Ybgg_m��i1��4-�jc����k��^���7Ë�xZ�A2\�E�>{p̹� ��XX}<ɧ��[��@�dz��֢A=N�V�ֶL�;�n�n���%R�+�T�ev�6
���@ãߝ�C��A���pB�����8K���r�Q���4"��÷&IJJ��R;��;Xh��Ql��������d��RP�*?.���d;T�|�����g�(�-R���ѻ%%%�I�PU��ieSL4���i�$@��J:ⵥ&�Z��]|`D��ZI��H`W��Y���3cp�B[H/-�e�n���ب7D+����ɿ����V��%^}�j+(�Q��G}l\\�|ي,�<�)s4�K�_G+�����̟>}�������я@�z�/�,��/��(ٟW�b��R�o��^�����%��|<���d��8F�۰�����z'�5e8}`V	��B���_K<D SAǢ����i���P�4�T�׹*ԭ��$3�ٌ��R������UHII���1r�ױbϻ��{Wﾣ��C+���.=Q����3�Y,�����
����%RILίm+G��3���i�N�Z��e;*J�RS-%eAԍOL$F��Ʀ�3�HjX3G��ztL�����zV���]o@fo+(I���nXDm}��F���Hϸ���և�YA�K����f��kH�� �=ۛ�{�D^U�)6���W��=ߠ������f�
A�KN�VT��A:��4Q�4�*wWix����R�t~}�~yZ�5�/���3��Ύ�v ��H�s�ټ뫖��бY�2����N��+��כD<��j�sq�d�E��m���O��Ɖ�}���e�����������*��l��h-~��ʿY*�*U�ojtl,Ubb"�m�ܷ�:u2���[p��^i/	�755�<�c�	Y�a䲚7���*I8_j�cxړϐgn=[��>VUJ�ʪ��%��_�D�O��'7�X0�3k��x�F�k��V0}��2Z�Hr�EU60�fҮW����w��Y�/2���m�~U��7,!.��H�m����׷��[�b=_���vM��r-A%A���/��/_�OG�R�۟8�:�!<H?���{݊�k26E�̑k�B��Ɗ$�C]�-�E�M�U˯\����� ```�)?�����uv)-)��cחԅ��]�ɺK����%2�,,�FCi� 3��������vg*
��<�]��MGCG�Y���Zڴ�Z~3�A�ۑ���8��sv�^�ׁD=�A,�j�??�d��o}���)�����
Y�.����5��32ކ�����Ȱ�Czu}��U�10(�k��0���[�(��&��2�Er�O=�%��y����ƧXu[��4+�	 ����e��&鬄IJI��ʌ����+!)	"WBJ*��U?��$��|~��)��k�svuu�SX(�eNE�/�NP�333��^_~K�G�p�����ϯ��'��k�a�ϟ�J�����y!Y��%`���H�Jҁ�s�Lϗ}\E̋�]����a�5J�����CS��A-�����JWX̧������}�9�TpS�@�������)֘�B�jV�pEY߿����� �~�?�z�u�<f�����r9`��@mP���z����v{��0������.�W�ű�'��|�D#�򝪡�F�n�f�?�������� �KK���&�2�h����V����)S$�&I���]�������1��96hwE�����NL������'��\k�	<����oK".~҈�OB��骪�l�Z�d��m̍���#"_+��O������J^��	^�� �q�)�A��?۝�]� ���L�~_1��ntn������iE�VT>r�]^��>�ܕ���,n�Z��_�5s9ee���xy$��gpSˬ�$H=eձp-!��Jf�m�Ro���6�z.��y�O�������	8r�����,W��F(��8�ه5���&�9ݙb,���Ӥ�K+���������!��k��	ГAQ���lz>�{�6@��Б�\=�&KH��T��b��z��L���;B�E�����f�zu�8���m~�WH���b�R�<��o������h���>HN�&��@j���:�4��=ۆ�3�����j@=���]n>�B=㺹�����У��Tsff&:::�Js͋����-����Dtyc�'��D\t}���o���C�E�냊N��
��(��y�9�@�����D��Vn���\E[�U__?��R:\��w0���x~��6iU�.;��\M�9+J���u����ȓ���f�e9J��Pp�UL�LS��u��@��I}����![	\����<��Щ��Rd�(R��@�?��H.@�tUth�I�QȕN�d�UeR||z��;�D)�8���܍ �Q���r�Ew�-���y�5������!AV9��XP8�i���Rj>o:�y�r!"ŵ�@I���6`U8~�vq�+�H����۷��	 ��x�N8��	�'����]'�����IK����Tu�W_W1�D}�*���7��ii�'.a�M�p=1I�N+��`8�
�7$ ��&⣣����B&A����@L);��h�]By-�"���9���9.Ꙝ��a�7@���}|�6bt�?�%]X�x��D#�����T3����/H�Ս�>��_*kcx������;�M�� H�3a5���>q֪�����":/Qb ʱ��6��A 8����,;��� $�cY>���P�է�~�M�fCC5�Wa m74߽�{��^P��fU/>���I{�>S�D!���g�#3�OOO�n>�D=�=t��#����{�u`���Wt.$zJ*��^w�y��J������-��^���up�������Q�W��,	}�Cm�����r�19<��1�DA��mvo�P(�R��&,M�dm��~ C��k�f�� /;wN�҈��///s70��ݣi�cs��q"z(���t�j�窙��]�g:��NSõQ�����jS��0�����	\fi�)μ�c����4���A�>�א��6B���Js��/�<� L䂞a�;L@@��O�������l`H���K�w��B�Rԁ�5H���oD'����R�Ce'��pK�ʪFC�R|���і~%%,3uvyѻW�rV��+*�99U$����5k����(OO�cTE\����t�E���vDy_k�AEEE׃TT�\`����v�v�88k�yiѦc�ix� �o�ӹ�	��<��H�}�*��?NnԂj�f���n�|?���<�	&tw�d3�nPH���h�{����	"f�H5.�����Z�ܛCFH����/�-�&����X�nH�#d�֟+�n�]�3���Y&W.���J���q����<�X�J�%�J"(����u[uo�/-U����v~7%B�6�]�+���$\��* ���
ڨ�|K]j�+�~Q�%%�����β�Y�4�������������ջ����%[����7p�_�\�y�KǄ`�y��Ck�[�T��u>�Vޓohh(i{���-����d!�M)�]%�{?Z��!�f8{��B�0��%:F���3��+��ho_-Խ)�B�7Y�����P�M��բ'�������"�d���j����#���733C�����CJ�>��
xldjV7��2ƶ@�:�YDt�{�)""�kU��t�-(/��JB��bl���0�&%-�j��!$$�5 ����OH��Q�ܚ�S������y	.�E�QeQ��`�e�L���b%�:��h�;:V����ψ'�H�t���J���maa2�$|����2=����}�ϕeNn�F9&nY9������WF��S�d}���`,Э�ihhX��:P���R�i���b���j�&nu1x�H�W������
&'0�}���J�n
������R?8�k�٤�4":�̤�#Ā�v�ǽ�8��h�N���.z��s��[f�6+(hj� �P������A��H�E������AsG�P�_X�=m%��r��U�n"��؜�N"91
�ᐐ����[�0���N��;�7����#� (��관R��j4�B������x ���h@1�� ���ݹW\�uTTT�A��%���3۟��NI)�TV�	D�pdD}�i��j��^=\!11��x&Hk��w�	+����pD$#�TB�~@`t�/��uN���� ,MBw1�7i�رyxh�T];:�t,���ՃVq�ޱ ���J����h_d��5��zjj#p�zH�/7f�{B^�5c���r���'9�x˟�G�"��
Q}�c8��)�b�DD2}��4��s�ON��TSSSw�l���=?�4��y[�Ԥ������@�0�e��T�)8Q\���o����L����s�\]��=�4s��C$@�of6aak��@=�%�w񦰏���Evw!F�� ?����'�\c1Q���uh��*�c���� ��2<cъ�%il�����W��ٙN���SWk���e�)����,`��Q��+��z�J��%��Q#Yb/�H�5G@�*��k�?$��$�f��stU�DSK�nO$M���dd6���F)]B#�Au)�D��hӞW%�G���D��>V+��X�� )��adbR=A�cҨ�����U�	�Xl��PI��eҪ�����..����C��$#����l��g` ��w��e����J�.tBS����P(Mq"L?�sڏ��׏��Җ�a!!��J���_��cz>V���/��� �dz��.���4�Y�Z:�|wׂ���!)��?��捲�y���	������0C毀�2@�I((D�	�����at�(��gQ(��Z_B��uSU�h�ү��(����yDwVQ�`/Wdnf�-�{�'
צ|��#��7;�q�g��H@@��S��~�V����$�7�gg� >#�ޗ����׉����@2�6�����3�q����U��,ҿZJ��-��ػ���2�t��-�h0;�Y��ք
��@u�9����xBULN\|<ëE


��ќ܍v����z4���ڛA�&䲹=짹�L+r�u
�eOsY'�<��*���QI���L'���j������aL┄������,ب�v�g�(y�c�|��g�_�x�ui��Nt%��x�u�"�6~�{}s�=��l@� 
�f�Y4���󂟛�U�x��#O��)��o�ʧ�$id���4no��]D�E6��'%}��W�|ʜ_X���
'������3E�ۑ��d���,��H� X6�쩨�$F���#��Zڙm$�#�~��ѧ��a�}3�	 J6��2m]]]A��Dooo�zwWW/���I������4���_
���-//��1�[
Չ�(/��l�Y/����(x���ʮ�R�|�պ���#
Xz��"���<)0˕	� ���dk,У��:�����a�G��6�O�O�y��F���P�5h�FA`�#�E�^_FGF>���������u��ӟ�-���_�� �z I��q����\��0g[�A��k�����𛛛���z�ړGS�U�k�N��M  ��᠏q���rs�xפw���f�w(��o4�DF$�0-��@��������"��zr1�.:�<���"A@r�ru����!�9'���p������?��&p�a���00B�v&�%�Ζ:2��`E��pޭ�O������+ji1��,v�}�?�?/p_D�]�}s~a���8 �R5�+����d&5����V�#��-�u��|1�FFF�<��Η*��?\P� ��h~�^�l����g�:�����x~��va)�b�M������[�w������W-/�a��Uښ�⭋(��T$�b��qػ��(}��#:8M]]�^�2T�7�|;::g�6��J��^�[�i&7��ǳF�n��-��||2}c�""���O�(�_��r�|�Ҵ���U}����Q�;6!�(z �<7�u�22a���3�y����~`\^��tk��4����Jչ-��n��W\Z:��x#9MSK�f��OH�S�?��;����אJh*�D�2C�lBee��Y�Pf�*{;�R�	YY�!�ؾ��������?���9��q=���x<�� U��Τ��� �_�yQ|��[��n��E�ѩ��c����;G�E|����1
�O&'�	֍[S���-��^��K!ıOu�%32�mH������ֳ��zb�����|u�U�۴�C~�s�i�W��"\wR�!����$(Ŧi`z�CRC#���r:�6��N���B�Y��r�$$%�r[�P�:���!�*�Q�WE/�u].�)+��i.�I=IEe�I~�z� ����1X��B��������?g|����p;e��'��sss&��2�ߖ+��D�d��}�ly����/p��م�5��8�?f��۾۶�R� l�rE<�ll�Yu
o�R����1 �YK ��Ժpܟ��є����t3c��u�K}���*�����{��a;�ݳ*::�f�WĘ��#-�.�'����O�9A����lw�E�� ��tJ�o.2���?q,mܨ�̓-]�+�Ș��ce �����&���TV�2�LL>u=׳ kTVR��?t�	�����U�!��hyh���"�wN��M9����wz�7�L��9�Ӓ��]�w;ߦ*��V�S��d\����k��߽{G-fv�ȔSJ��?��/��	<�H&���Tʨ����>���^��dVp�ΰ�߼���==��q*���7J FS�w4]г�P���:��dc�����n���U������/��x��U��[����(����ۀs:!]��۫���~�wD��N�N�U�m�F��������[�h``�ֿ��MꉐeRaa�}8*����i���&$Piz����`+Q�C�؃z/H�
ե�$��>�9��=y�s&Q���~~!ψORF�/�;���<ʽ�kUe� `z�7g&��(@���&��F�߿�hHN�N|5�z���i#��z�l�2�I={�=��?��S=�E_R8�Uv��+"
0.�ŗ���~���a��M���� ?��[�� 8�X��/�����{�0T ���&�84��^?��OD��@H��T s���_?�bbb�:t����+i�������z���������d#W�
��i��}gvB�5���(��_������RH&��J|�t�o�U�2=�Y����ׯ�Y7��H���9o�+�K�ٗ);��IS�5o���S�v�X���3��������;���1e]���>-^�9�WQ��I��hMGHe�T��i��w*�**$Z����Ya. `<�e��}t�<�N��L��� �[�y���e�@u>>>�)�FY�oT"��߾���W�m�5�ݕr���1���%=F�o�5x�loo_Z�s�ō�:p�Lb��Sy��}���T�_2����>����������ֽ�� ;@<`������Jg��IX�\r��:gDIpE�۷oՙ�"Q� ���6�/_�T��e�����j�MN�s�Kҥ�,���Yxn�/��zF^<66V�.}���ȏ��T�pK_j)�# ���|��XK��?��'��r���"g��+k{ݗ�g�_/��6��#K�iii���g Q�XX\b�a�7}�ŕEթ��OR����ozzt�M!@�O��K�B@P���Z�-�;q���$�ɫ�.��Uq_32�7� ���H��Vҷ��'��������`���H�?c�O �|n�W�k{H&^�z��E��_.JD�u�걠5�ʳj�q&}�������L&11�`^�j��?nnn�/O�R�XZrj:G�Y�݇j�	��{���­�?-��(��x�]E�TXĝI�����IHH��Q" '3��ćP�PYS�>���֗F(~��߉	Ki)��EB���:��poH���Ib�W,��C��22>F^^���fmK*�r�-����.R
hk�4�J�Y��r�GV���q�Y�vAK&��{�j������.pp����m&��sڸ5�^{;���_����`tw�5�'��U?(\wGG�
#���L��*�#3kM��>�ؾ�c���Y���-�:LݭCD������=�{�%E���4�\s�:ݴ?R	��r�E=5�|��5�9�EP��6u����~�ͶE �?��������T�+�4�͛h {�*j?q[��5������BPgD�ʋ�p�?�Ro�@����яJWB��j����RvaS�bx0�YG�mRo�+ئ���H�J�+�,	���x���F���b��Q�͋��e��r����c�&�DsbbHL�Ϋ�����.�+�����_��8�B�,�1���I����Ǳ��E;��,��^P�Y�ʾ�\��P�s��!�,��F�[J�K���D��'�]])t��FF�֟�pq)��6�@N\�����w�`�R��Z�Lbb��v}%�o�0!�T���N�Q"����3/_��7040��� �p�s9N��_36���ʵ�u�mo]xs����"M�ć���+��U�.�,�F��-��~=,X��JsO�V�奕3�?���LDI��w�Ni+�q������K��Md�k���u�F�â֘�M�,��"��P'��� ��i�I�=[R��{`u������`��ش�o�X^
��/.1\T{?�RS[��ի;�����^Ն]�N\i���toA�G�v��������x�O=����5e�nljB�U[��:ZZ�<����C�ᒞg^<x� 6>xdQm��zff�͐;L��>�.��ߌ�u�--juMu޼9s�ȑƞ����@~�+��M5m������CAͿp�����gQK�4�"~��wK���Óe���9�:���2���y��*�-������l�o���l�<,��X.\P����s01)	����w/�lƱ	K.M\�������i�L�fe5���1��]ʾs��k��
�����.?՞�n}�"h�����_�I�?T�]�А�l�_0�V7/;��P}T�r~kc����=ׯ_�qs+���w^d�@WkQ0�G0�Ccm�k��-Y��M(V�:�5���`��W9��4��'�ni��z��])��N{#���7:�������f6�ϩe��cf]�U����y��#ͅ�����,T�^;�&-)IwP�����kӃ5���"��g�^TY<v^��&�`󰖛�Zz7�5�F�y���v�@�3]XPO�_�� �8���s�_�m�JP]?�:��Q��m���|�g8�({�]����qG�I�\�-begFh/o�R��lV��{߱��_��w�� ��t�<'�015�����C���c���1����Iw]��7~{�L<�ϠKԢ��j̙��&�K}�ұ���cTt�?~�^�)}�'���^Q�r�� Ƌ��W���I�<&����l9��'��4��98J,kL��Cid��}�mIs�>������z��UW�X�[��[�\��0 3�˰�T
��4p��4!~�{���ӽd�h��T�=������宗�0>�,wǮ�VM-�"ϯZ��m�Ai."����\o���a���̸������遪���^^�~���}��BsWd��\�UI�
���W���NRh�^M��I(�E�4��m���[�б,������YJRj����&׼����g��&�0_wIX��ֶpط���_�~��J������~c���B|tH�,8�ͪ̕`�K���!{Ҥ)u2\�}T���^^���͆�S�^�7�+��<��v	d�Z�kd���d\L������b�;��8��:��Z��.O�p���u%����:���8���G��嶜�����9|BBZ:.S�n���g�|}\JʸoE�9���B0𷚕���������\��:WJS��oF_�__Q�<ޑ'����w�F�r� ��'>/��i^�Dp�-C_YW�CCCCPu@�ˤ��� �m	��k�����L63��h�9SUU�j-��3Q
5s#}y��������˵?~�E�ZZv����h��%{�P��ZOɑK�]��*��1�Wݴꨕ5,a5K�bfb���_9T�F��v��ٌ?������ O[�Y�3�~��%�k99�UðW�� ͪ��)���n���d.�cP���;w�(߼ip/��Qx����Ø��,*�X����"#-\��V��f��5�r���K� �P��C����{�/�hZc#��sr��ZGld����C,hlm=o���������ч���2�-����̖�{��,�O���g����q����))+�4~j���}>#�;z옾��:0{iJJJ����+�X.Tȴ����^;<# @�4<���^Wx8��e.~~��勘Qw;�z[5==}����ϥ�]111����A!!T���){����Ћ�k+ν_7�K�Z���=�t�@�Ǖ�Y��gt�������q�'N���I�X\�.o���Cv�M�|�;��<666���T������}8 \MT�i9v㚆�j� �p>�`\Ѥ��tMu� *�j�/����,���O�m3��_�~Uz��D�QY�}�����#M�?���*$2��#����#:`���((��JE �Q����/6.NZS3�nɸ���^]Ʊ8��H�����sJ�B~����~.g�S������ם{~Lt�:vu䘅���T2��|��?z�(�[��I���c?��S;��g&�eT�Z�hWx�K��G�z�4`'���(��e[$VHXk��W�<e�qzɅ�Hk��
9��k�A)�%:���J�틋��c��؞���U�n6w�<��Me��~�*ЀC������8����Rw�DK�v�n4C�8�6��I��6�U�:k����0���F�D5


�7o�w�M9z�سg��n~� '�X ��wO]�l+�Os��}�F�͈?��ys������2vsc�c����h���Q.���^+�V�*ڻY-˟�L+��*>O����Y�s�xu�k�:��,Tڎ������k�o�yYa�X�G�����J��[T��v��Ԫ��aU�#b���ľ��%����sk��� ��j��M����r6Ϣ#����-"��������3������d�Ot������ ��B�!�j�jPX�S�(��fL=F��3�7C��$kp���kihm}#׼�C�Stlj���N��R�JikGP_v�aK��AduF8� �����1�6vv��Ƣ��T�C��~����/{qoߞ�3��%%��(�T392�F�P�`^GJ�K��.y���(+=	�����<+�`+[�Z�V�ɬ%�ٳ���Dv���#\)�^����\Ct}wZ+:g2��S�� `_�����|M�ݻ���|���BL�'������n���_'U��Pǩ���<>pEi�K��\�w;99 kI�����(���������O����%HQ�>{��m�W������?����G	��F�."R9�3F�	j������@���D�&�t5��Oް���3�����x����'����$|i�YE����#����@��q;fV֛�$���O��Z�����5��\2kMJ��Kd/�A�k�ƒ�-T�����Xnv6"\6����=q��ƦPAK_��˵�)��0u�k��I�4��K��Uƃ� �׿���Y(+�JI��ʮ�&_`�C�����<��~��5o{�#z���m���W������z//���긋�^��&!%�`1��gy4+�~U4�j�4���� u���H�`��V�Ee�]�U>���}�)
��PơP&�oci%�O�<3d\]]���]kL��'p���zS����3� !��=}���$`;8���nl�zmuYucM	:��L��)X�=��n���}��S����L5�.�<||,5d� b����6����Y�P��Nti��;!;97&%��.�ɢ��=�
 v0��	^!�̕�::��̖����ۯ|�v�<�vG���s��k�����y��j

	��@:͔�;:�F_�6�-��y�QW�mImz(�
�Q��}Jb��}�Я�N�za5��{5ڥ��c��n�}�̈́��`�WƎG��,���#�in��#4��������R�V0��e2�K��3��ebf��OCNnWs}���aee/��\*2��آ"m���V�r��M�u
��6N�̶̨����&~��Rbbbj�(��	T�{B��'��>��2�N�XER��c��S��Ԕ�Πՙ5rrr��Q�γ7�F1;�~J�MJ���
T�(���Ww w�i㛐J��8	��Sv��<zcfa�pf?A퉍��iT�hZ=-VWZ�ȼ-�����Fh�y�;=J.<xP.��hd�e�C��<����v�st�^��'TR���#;;,�pH��41���qT~Z�L�]5�1ޒe�#�8]uu��2W_���Q�0w�(y�W�}��>7z��DY��:��@`L*��:i+X"��--j*���}
ge�x/]���>�����H#��C�y�����'v�[h�R�&<����+�r�̫����?w�f��0�+��I�c�a�A��bccQ���l0k�
�;� 9�fG��h�U�Bvɵ��ˣ�t�N٨b-�F>HJ'�Ϋ���X48/�\�����$$$�uVn*:N#q�W�� �Cg�x$Nu���jv�}��G��,\궶9�dس�Y�X���Q��I��a����|�#�(�;\5 �i h�n�'d���F���T	M�E7 ʹ����C���nc���R�] ����N���K{�Ẍ�e>���7��Vnj:(���������\�\k�. �ƙ��俣='7zt�j�=��|h%$$P/+]�1OҪ�z������O��m�mЊ/���'��(ϧ_ �t>ҡ/ߌ0]0f"6�����
���8�ۀ�/��R���p_+D�Д���z�P�9 �E`��9�`��Weu����_�~��NH;.�$��P��ǻ���������³�ؕ1��_4���AtX�5٣�}��U���K_������dڻ�2p5�"��*�����#�������ޞVIPP��`XWWw�瞱�YK�R��������ႮT�߹�cAu�ȹ�-��3� 䢤�4�#,'*r8�ͨ��Y���0�eH�)�,��IC��Tpֶ66����9
�}�����?��N�����*)0�L�ˋ����Dd�75Q�.jĚn�Z�	�6��n�"�jdQ�Ռ*�����m�F[d���W�����EP���t�Rs��"�×�Øwb�@�р���^��n �{�������?���Ӏ�J*��4e�d�Oꀿx�6�D�[�,N��m\��$y:�������\��o#�G40`�4���V�El^�:j�'P��Dʣ�O�7�E����X{tt���T'�Bd �*Wq=���?�P_��CGtM�����j���ղ����D�$����d�R�l�v9�Nȓ��2�m�:�z8�S����7d �QVwQ�.'����A�L�
��N5-�p@d�A�5@A� �˅�]|�M+:˂�93h�o޼Y��L䣍1�������~�(�'��j�9�������ݥ�x�E2���Aջԛ����╀,�/�"��vxf� �tt�����Ɉ�
�ٍ�*�#����ظ�+�vzD�]S�MI��;~%��h�d�(Dט�2ס�P�с�w9}
�r�HS���r���$��'>�����0x���U)�����+7P�)؂@�q:������;,�	b��҆zɫ�R��)��Ǜ	QcD���˖7�����Uâ(�/''���2ps7)��ADJLJ2���`�ߝ�����b��.,8�
٧"���Y�O,,�`��� §�{��(���ruJ�~N
�����7���؀~��B
	m����
�~�K hp=�F�;�M�Gt�*���������cdD9`�/^H��D6��;�������Ld³�����;�!캔M-h#��&����R����p����=�U�]|����3(A�~Htn.���|2:$@!B�q�>*`i�aXbA�ڂ��gJ�v�=�}c�/��'o�H�m�� ��vR_rz/�*B�]��c����Ҕ�R[[�ތ���:phȨ=�*
� 'O��{}.��7G�4�H�ZZ���p�|���/_&�T�r#
X�Kߜ�jH�������li^����b\�܆����딢n��礗ѯ�*��?z���~G�ӓ�ϊ=788|�:-1QyԜ�u1�����2aM�E��O==�ƿ�t�+$�4Q�t�C[�*P������*�R�͌�=�lUUU2�i]-Eyy!3l_�fg+���6z5�s���ϟ{�,#��h�o�)CV"Z
��>1��3}��l�9F�Wv(�{s/���K�8�<:�ݑ����n����~g���.�Q��AC M(�_~�4x�عʯ/����F�
ߠ������� F®�K���,���f��
�Nͻ�|�~�ɍԏV�TƗ6,<%Z��uq2��虘����e�����������aQ�-3��h�/ou�~k����U�
���Ӈ؟x{�1��z�/����sѯ~ 7�GԀ��]�`���<��� "��l���*��Ap���?�@@ښ�j�MAW#�	���k+�(�x��F�s��Ͽr
u؅�[_uu-b�W������Z٢hWvũS�]��7wEܻ
f���ăv���&� �f5tBQm�3β��9o�K/�����\�b�qth���R{��)d:͙6�M9\F�D�e៼;��#g222��<yf�2}HZ?5�b���9�"� B+�4�1����:���<id���ړT\y���%%�^	��r�;��n��⽸�DVo��� �eHY�اϞuM]c!SYt�����LZ�hogՠ�O�!;'GZK��m�UPPB��3�#�	��+Q�+0�wOJ�ݽ'�%p~:�IKKl(zWʾ}���\���E�����!0$i9��撒�ռ�qu]2	���%;]�[2Y��f�l'g�4g�����M]�ȩ�@S�dkKqC�[]S�G�ܙ3WѾEʛu���+S_�AV�A�Sb_Q�$� �eYg��X��h�Ց�9�#/6�)^K��q99�0jՐ�H���mf=T�p<A!BY����!�K��O섧��,MuTU�>m���(E����ߨ��-HZ��r���Γ}����6�O���?��ŬC�B!�D"A��0���=�ɍ<���G�Ӕ	�|`eq&~p�Qk�8-|#�@s��u��K��{�cm.�|��&���ƣ �!8��paJ�N��gf]��5���#_��5�j��b�;�u��Ϧ�ڃ�y�䉠���<fTf��nl=,O�������>@��?�F��5Ͼ���Q�6��/��|��#;91�%��Wz� ����{�"�T���6?�y�1���D.6⍯�����+̗lh��G&�
���g�?�9t-5��1--�L�
�M�� t�T��gi���e���`�߽O�y��VY����yӥ0�L�?u����XZ��������k;zSZ^��x�x��s�@r�᫬;��3MOSS�
�ֻ���y��7$9t�%6q�|���u� 8A����l����j�&�θ��n�T�DP���xCW7*����GA�>D�����u?��h��s-:�4�7�~dr��X��ݻ<4��o�+���H����&��� �Zh��� �����~����_Q���Ky������V��+W�E�F���W�'��)�{�|�u���2��.d>1�IP*|�s��f/^cc�\]W�I����y�	�e�"����BK2��yw9����`6�KY�g7��ۜs�6EB2��
K"��$-Fy���t�˓%=��+f��"�����&|E������[�5��
'F΂��ܴ"�����P�T�H;M�ay�C�JD�&��2z�����~�7��S�A}��+z���܊ѡ!+b���g�N����W8�n�+�|o���+`{�ۺI��N�@��q"h�����qB��|G���f�g9-��@��d��"��Zl��e���a"���<#>��m#D`������x��c0� �^щ�վ=pN�hx]|���L�z-'=^*��9�D�6��5��#�w�R�+�R��\���$4
�R6�
�v��I�KN<������{�����
rپ�'�#��G��f�A��cK"�k��&�6N"�Q?��mλ�x�B|~��R�`Y(d���`�~�Pp�i��_��ZH�����G�<����]iD�j?�ٳ(��}}wz�^���%^��GKA�I�q��J�ߧ��ʪ������	l$�&o�D�{큼�m˃�%���zԴ�Us����'�Cr�%�:���J]I�G�J悋Hs��k�w�}����i���v�����XKJ *z���x�|��v=�>-#��v����x�q׼3��
XSS앟*D�D^����}$�t��y����_����.<�x�����n�u�F�S[6��yo�ޕeܲ:�A$Fla,�2i?ޓ_�#-���Z2&<�n'�3V"_�+\�ڊ7\)-�gQkS&�|���'��PU)��[���<f�8����+g�S0Ba��|S6������5��$�A�b�O	���w��<u������t��u�fD}]o�덚�"q��{�w��d�$�IB/	��v[�L����z�!J���/짹����؏�k���n�=�s^nƪ��eE=��R�7="��ĥ�X�\��*���]�Չ{\B<�w+�Hd�LNN���g���ّ���z7^����_�X�}���2���P����7�@PŠB�a�u7�K�u��N�p?]�^b�(_O�����8͔ܯ�'�۳	q
	6ŭc�2ý�α�x�P߯O*%%t�#]����������5��<��]�p�]���Ox��;���/���SӖ��ق�ۺ_���#sN�^*��G=
<6PE����8�o!�g�[�Z�DA��Q�����9�r	M��^w��Trm��.t.�ki��P�\��j��Z�jKީrr|CZ�j7�ͽZGoh>���0I�F�f�)>O3���A��.�x�-;-���JŒ���x�����1��[^��޺�j��5��\��	��NTX��z%K�Y�ua������X1|�u�B�ֶ�<����Q@�j	��nYס��{{v�x�����ۮ�¬O�\W:.�H���-��
��Kwh_h��E)jBK�0{j���vj|�̏i77�	�oa蹳�*���^-��YId� �:��c�|��D������"�a��-��֎��&�%���j���Q�'=*�`��!�Ԯ%��$Ba;&M����]t��x{z�4h�@�o�Z'5W2ț�~`�Y���Ч�ֱĄ��!?���\ ��P8?�����W���	�B������5��*�n%Q��_8����PH�%В 9<);=₷'��.��m�MС�wt�B�/h����΍��_�W��0VOW*v}'��mW���x"E�Eş�|�t;h��:iV�s������OW͝�> �a��ӣ(�36�Ÿc2]��]��.�9e3���8+���Ლ��~��$Ey����]++��o��-�CP�n��A�Y2��&�t\��Q�l��2��.�1����v�C2�|����D\�GO���k��j�W��|x|uk���]�.�'� �����"�tZ���.�.��Y� ~�
��xv��W[|�x�H�c��pd�~��o_�P�S��U�<�>���C�i�4L��咨ӫ��������far}m�_����X�5!.�d���\������@�Sg�5������7�����̲z�3��s���P�����hz<�O�,|s�>&BwX��U{,����X1��_�EfB1����2EP��v�s����\$A���s88�eɷsX\�1�������k]���y{�:}e�9OF��յ�RH�*�S�/d|���X�LD��IS�=�S>vȳ��v��d��yfd�0��[����S���,y')i��µwh+S�
��2�$v��Wv��\�l��]�<��u�)��o{�ҏϷɨ�q{c�F\��Gl���sN���Yk0Sw�	ٳ������T��my�L�,������_C��,�ȩCw���C��r���>bC	AΩHǦ�����P�o�Zʚz���Q=ى��~�����������"f��+ ����p�i����tI�Z�u>����Мs��N����*s��Z�6���ZB{�C����Cf��u���$�('v�����'5��~O��'M��\r�)xE������k�֦x���sIO}�Z'�(��>�8s��L�;YNڷ����|��)@��ǮǼa���{ܮ�qG��n�Q;�Cީ8�П�r�_��_��.-���2	�-�Qt[�l�ۿm���ދ�1쭴E]u�����
O�L�yڶ����P��Į@�w���N�8P�9���zOxk߉�t�_����FU�n#uXyy���1�*{��b�6�{M�x�ެ>��1�����
�_�q�	�s*�B�&cz�;q�I��'����Ho,��PX��s�����t�Zct�ڂ/�Y�;))�UX�(%&V����a�~�e���B�ֵL����=Nz5����JX�2:<�R�V����hZV�ey>���K��n{�t�/�ZYM�u�6��܎����p|� Z��c3ZY���O_|�>�c��\�p�Q��a���*��k�}64�/^�}»G����C�4�nw�����>��Mkf��1���la,�1O� 9��g��U��F�V����=������x�*�gnZe�:,ƙu�6�$�}��I`�촯��]K̊��1jI��y��J��O0��1�3c`Z�v�;�Y"ߺ�3�Uf�_�e4R��8O1D�툹��NE��N-Y��l^	��˄���{��p1���߿������~�a�,,)�:pӠC�o0�Q_���\�3�|9%c��P���9�w�B��H��u4';��qvv���	�"M�qxt����4`�c��"�����r�#�z��; P�g`#c���w�4�k��ou�G�	 l+�⣑�������eE�u�Z1ۗxbyy�5�� 櫇����~m���?�0�iV�DwD���#q���#�J� 6����S�*J������7�'ژ��wk�\9�Ƃ�9�X�X�������<�H��9��&����잝|tb���Z{t���2޺,]~�3ֽk�$��d@H3E�9�d��u�,!�ŋvs5�mW�/"��N�*��3^57��/{΍�	��p֭���ʊ�N�6µ��Y�3W�fn�N�]�k�.!�$��'ꌸ��c d3ͥ��h�|5o`��	�H �]����T�C+;JT���fwp����@���Nh)��!߽h��9)qD���m����~RX�=�8q	����ó�W���\�7i��W��mrN�hSS��c
^Ẁj-���)�����+y�z8wmhž���V9���W-vZ]x\��|a ��L�Dgҙ�L�Np���̴��{}�@�`���X�/��2���,���r���~µ�umCXe�H�����Na�8��}H��\v�t#�<0�Z��д�Q�ڞ��zM6uc��	qu��>��[�"�U%!�9Ղ]�FlLVQۚ���b�E+��*�L��mm�I��Ps�(}�鴚��v�t��~�|�o��Ǡ�W���{���	��}̐�R"�����փ+M�X>���j����^6Rއs_�%�f�G-}��Zm�J�G
����KZr�1!���n��l�����������ǳc�27�eF��da��~���]�H�(�1iW��k}�0t��zkPjߒ���>K:"�t�*KJ�A�;���N�bWWW �����>�͍%���qo�[z�q�����7�٢w:��D�`�2=9}h�@Ȗ�ni��L�۶��ox9���<rD���z�φ��<�X��_�8���f������Z]vb�0y��ۼDӚxs�iɲU�}�	�d*�s��Ic*��/m��Qʝ�'��x����8kV�Qʦ����3O��`^�v:?���*>,D6�s�?uN�	��3�G�������ϻ8��)��&��[oӳTw�q��2��r��	�I�^S�s����K ��!�j�Jxdk��9��\b����15h]e���N���@�J�]����ͨ}Q��/]��w�����e#�3bfS�ϊ�bs�t+��x����5�>���P�g�q`ZŢH�mң^Qa�S
6�u*J��^o6��hً�]�Ou⃛j�0a��Q��'�B\B8�d~۞��v�1cs)elAnt���~O�D�p�����Aj��2��7�x���r]���k��%�������5WD|7��������L<�9�u�C���,��?���|� e��P�:�6�7�
���"�ܻgvd\/KS��</���/1k��#�h�Ԅ��u��_�zy�NX�˰l�,WG�@4X]]�)�n�0nPҰu��������};�lnط� �@46����KN�WK�����n|Z���Z��4��ey�k�����%�|�6B�W(�z��I�s��~�6�N��p�qSc��m��+����U,�z�,EJ.�ZD�Xj�=�S O����o�v H�Gu=��^�O�Hۣ�}+2׋R����~���n���T4a��N~`p�����@�z��D}=����P���9.��<Y$�"�>r ����*	
)jB-�[+��,g,�6���`P�8�?9�9哝T>ߕՋ�r~kr`Ҳ����I;V�*��3\�����E2�6��������T]ӥ�ݮA�c����:Rv>��ZVH�t�F�Dn����e�H���Mh�..�p�rx7��N/]�0�|a��@�������������:��U	/�90Z֊|`J�k[+q��r�G�4�Ӱ���	xϻ����znY�hR�w�P[��O'�d�f�ԶeX����=��~��9�g����B��9���m
���#�����e�7��s��7昼䱼��6Msp�qN�L������Y\ ��#p%��Q��%_p>V��O�+�@��?p��'u�m<�96ȪrT��,�_��ʬrV{m�Ј`�B�NZ�Ÿ�����I{��KB��2�J�u@&�>hR
q����	q����8ֈ�1���m�����_��Y�$Ľ�9CvLy'ѓ���rys�[�s��ϗ�F��1���s��k��m�+P%jcH�������ez�%��W��^�(���'G�g�Vߑ�ƃ�9_g�T��l]��L�|ڈZG-\P:�R�9�)��[A������L��z���&o����F2��Pp����[1�W��Q�4�)����_�*2$��I^&�f���Ϡ0:�b��q����h.��ةnS��w_s��z��e�C'X�b,.��u�%z+J�Z�E$\�'%#����ms�楡A���j��?,~�~0+%.����d6��Jj	qv6��9K�nr	Ml���}��乬���xI�&ٽ�e:J��m"~S��������Vrv�����R�:�����y�H�Q�(��?�?
��z���pWY�(��I���5&�Js�A����/���V|~_[�8J��9���n���Jg���a���[>�3��䢷�.BP
�D�9���Ɔ!���.��n�� ��f;�p�R�h��<���[�Rd,�qTJE����Iu�>u�nM[�H%nz͞��"L�E�ؠ,��'T.��C+JՊ-�
������\�`���Oh���"���łh⏲K���	qn�9"��m5���z7�;3�mV��2{=��u"cc{�6���[���]��Hq�'��� �����[��6 ĊI��{zz��}@TQ-Ip�N���xqO�	r��P�tt���k�zƕ�Z�eS-=.@LT��S���=�UT����j6�L^�"����Z�+����.�>��-v�;	��𓩥���s�Iq9��d���߸�sp�nç�����M�"�c?.񆙤F�oN����]U�ܲ޶�~';J�SX�R�8��YO$���1F����uX���s3z�34+��L�=��	���1�=�E=�ea끏�X���?Sѹcç�q�lE^��s�)K�2�8ۂ�!���C�ݒ�e�1��zi�#�Ld*:e�E'$��p��@t��J����[��8e@>�a����z�Sg��^��\P��u����x���\����T��+�%�Ȝ׶L���G���Ԥ����Qda�����iI��T�������^�k�͉����7ƴ���T�����-��w]��n`�o�:9=t����1qʁP%))�ֱo`���9���ͦ��r]��u�����|�_c���,�^��	�I��Ʉgo4��h���󹕧�W|_ ��֎2ɝ�@C��&����'&�OLX�����TԖ�t�2��!K�o��U�͔j#	ӱ�tI	�f�0�Z�k3ڦt8��\ה����ncyn,k}k_>�˂SR:~��/@$���\�!�K
���Ӣ�~��}l�%K�oy���W�W�=$xd�l�E�ذ֋~)���9�B��0��h�g:�?`�q.I�����予�{Ii
x^@Q2B?l,��3�b�I�g�����XR& 8|���]�͋U�O;i]��������\/_<6�61��^�f�2����,۫�'����s�N���U:����el��Kk��?O�w�����AS����S�����O+ ������籬�Y�#�}K�0��,P����OO���+E�3Ru�{��O�s�ñJ6���퇦�'���S�Ñ��Pl���G������I�Hu�⺦�K�kL�.��Ңm�������|��p�í{���Fj���H����')>��%I��[eE��<�/ �; �///�O�C��\���s�\-�.��Cr�1�g@�/�|p�i=J�X�Q�����v+���s���z	A����o%�CE�����0�6�����W�P��J߲�>Z���W�B�1i	(Σ$�D����Xݾ"�w�n�S�&"х��j�be�CfB\-�GeE��Oc��\�K�g�^ק�6��J���R�L��l�0y������s�6�;e�Z��m��F��.x��"���F�ǳa��ʹ�l|�*��\;�[� 2�i��d� Q��iSy����I�ʲm ��v<gtpb��Z�h_Ѥ�U�E�4U+g0��V�}�*+z�z�@�HĤ�q�L�d���W7��fe��+.c����	q���&�{�ܗ�ܩ$�n��|Huh�f�0�p��?���	[�,�PF��n���+j�Wj{ `�d���:�R
�;��7�ӻ��}B^?M�t__�Zj-��4cҿ��j2�yi����(M��b/F,��c�M@�����Y���uN�7?+n�F _����O�7+�c��r�SB%3BSݸb> �����a�)�=�M�o~?9�y'�|��\��ʐ՚Q�뤷e��-C�#g#�h��>��r�����èl1��~�I�PӕŨu���J�(��/�Ifh�>�ϒAE@aY#���6��f����32�Q�?��GR�ן�a�]0���6+��3Q8��:ߑ�[������ ��MJ�ŉ��$S�d��wV<<�>�p.�����ML�L���}����L$��a�a�}�}ɿ���1/����zzD[\�U��o���儀�4��"�^&�X޿�AB�� ��b����w����|u~e��ly��B	�c����M����;�N��:Q>��{یл��_��i� ���?�c�^li{�7�c�hr�&/����^s�7���������rC��W�M���3
i�4X��1-�N�� ��Ov�s�w��<X���( �,gZ1"ܾ0��d�YV�U=T��(_��z����ۆ��S��I���
 	�Yu�j�]���q�u�&��A��V���x�����;�9������țo�F��;3ހ���� T������T���J.F�88Qz�	�Q�hMT~a��N+�5���oee��4W͗s�����;J[<�_A#=�⽴=HA�&#I7;Ԛ�di�8=�n���s%�}�V����q���ێsN�G���N
�I
Z�G���3�*��Fi��Ɛb��o�'&���"y1�z�q����z���\�Ҽ��W�#��j�s�St�S�3G�����;�h ��a<�+�1�A�,���޺+}�&ʈu����R뮎��8����P�R�LW��.�ř��H-��5�\�N��]t��_�����:��=2�<�Ҡf���:&��7�Kq�^y��F9י�CE�4���m����/#��|��HD��8g��hF���$iӌn�^�i�.[�¾io�jQ6��pڹ��U\O��6/M�1��pu��� (������5�����{o���;mN{"d��Y�C�,�Ȓ=D(d�`,�S��첕5I��e,�2�Hv����`���7e��{�}�|���u����u_��z��{�,�cg��S'�fg�f�I�����30�WP�IOx�ǃ���k��z@G��"z��?7�L�-�B#�0*&k�DJ��t���v�|����=���V-գ�l=R'�h����7�����á[+��ƕ#!�÷�=��k��壺�p%o W�]���IN���D�N��n�{�lMBA���:�^u�������g�Z{���X�����:c���,� ����\y�I	���χ���U9�� $ �Bx�U���`{�t�#z�cYy��G���Je�[�n��g��,��*�9RU�2�i�Њ��[���C5k��#�fLкn��;Mߍj�/0��pn:t���6�l:��yKq~MU��F9���u���&mN%��fn����6U���7�Cseu��a4}��̀ùa��������<Ӝ�0����f!�svMǘ��c+��d���-.�I�eyќ ��ˢ�pk�aO�˽8BN*#x���[����>3]v
����<N���� (��������`��d��G�(�xi��i^ʀ�0�@�<���r;�+.q��L�ҐT�W��}�8�T:�W�ѫxѺ�И�S���Mo�aR��n&4��*�Lw��Ob���;�I��z�왹W��3�ND�2�,í�=0���	���9ߺ*�W�6��a(�c�
b�}��~��Gn���;b�}���A;����� v��������:v���.������1���Ď/�
�+{�4�$6J�Yl��ОI�p�"p���Ft��t�3|�2́�7b�ȸ���yod<u��&����q!�V9�59sj(l<m�e�tF�l��lI�5�m�Zo�fߣAl�WL��)حz��ϧ�>��'�(L*�}L�����i�q�2@���������?"������P؛8�\��� �k ���*_������q�Us���ה����o@�&�Y�w�v�򤡉;���K��*5���=bV�2S��<j��=A@u�}J��B5��HGUQb��ytZ����W�d�P,P�Y!��օ�T� �� #�5}�\m�m$��:f63(sJ��o����D:]�����5(w��u[�q��^H�٘p��vW��s�����
� �t�ɣ��c�������պ�W��Fj���؞ݏD�A�v�:l=G|���c���� ;��b�c]��0t��E�Ƒ�~�\��������E�x��w�=Ip����?���'���v�a�qaa�DS�l��k7�=���sȉzH��C�g��8�d4v܇l��(_;�J�5/4c�QJ��se2\AK��������h=*<K]�&�R�sGд���!�h�(�x��tZ'��g�����%q|�?��9h5���v�6�e5ol��b����,���y���W��S�5�nf��˥G7�:�u�y"���g��������zO�9�o���y$��/����۵J�M��D��wI'�>e�/��4�x�_��c�{h�b?G՞v_o#���p�-��+5�?e+���\X�Dy-'	�$����+��#����̟s�=��eE�|QQ s?��UՐE�P��;:�lu�<!wWS^�����m�o�G~�*���B����0C��17�o���<g�� �إf���qAx�\�?�g�0x�O�Z3��c���~h��wM��.WK����!���ھ����.�<�t�#��d���ܽ�{�}�)��z����KG�д�l6*��B�d�'J�)j���k4/��br��1V�;ހ�c6Fb,��f�P|��}�Z���]�6J�ֻ^0� ����J�Ll|�5������H3Q��\��1�>s�Hhw$
Q���6�uw�
�H5����.�9��A��|�Bp%y��:��"�#8��=+9��q#��"��K�"�MO����h̛t��Dl��l�Z�y�H����9��ͅ���ê�B�]3��c��~��&@� �C��i�L(��b���F�I٩gC�_
�Nq9X͹��_�*O�Mn�zI�17,^�!��B]S�lk���7\�������cG+y"�L��$���y�	JcT�|b�C��M���+̘3�cr��T�qr2�0�BPPP�j���mFp�Ln�m�R��	�+��ݜO��ZYM��(�̔�h�!}��g�^�{O|ѻ�V�$/C�e�l�I��Pt���S����?�8[F��H��ϋR_�����[�6�<4Z�`|X�h�u�AX�	Uˠ����,�4d���Ox����Za?��uB��x�˪�����ǩ�I�.R	�:��<(���/%1�!���������+ۧOW1�O\��^��H2o�2�N֩H��EEE@!�O�>%FN!��U�����i���b�-��Uth����b�{C�[��diDY�J�;/���ӑn������q�m��/Ck�&zФ��\)����u��#���[M��aI2N���tt[��[�#&��=8�TȌ��!��X'�`cr��B�Apvv6�1?��ݶ秀�lk̭hWF�]�;0]7�5d�iE�uc�W�xF�� �s��m�m�\4�Δ��I���H3��K?�
�����>$� み>UU��E��\��0�w�އ��y����϶�h�U�Q�Y�҃����=�w�NJ�����$#e���=ȗ�Ru��VHQ����k�q2di��'��ɸ��.� �LdW�6~,��N(�e	����;�>+K�"��}o)�E�.�l�����d>͖�b����������A�+q8Thp���<@Ë��Eu�
���z������/{�Nl-���E���P͝"7�*M�gr+*=G�9�uf\'�3DM�]�i�_K�S,�ty=u�ô5�S���_d��>���y��8�����ētt
�e�!C��M��#��x��js�7M�
g��6�d�'��D�T�3а�N!['� ;ʣ�рL+t��/8!!�9x�O��'=����)�q�0I���R�H��~М�g�$7ֈz&&������π��(a��$}YYY�<I��2]̙'h�y7TK`V��=@&����P� ��gM�Z�	tM��j�����%�°�k�:@ށ�1]3
��զ�z0�~ ���pŘk��ݗ�������_���I�8 r�r&�[2\������װ���	�=0�;Sd��ה�X4,Y�HsE�ϊ��sn�	�������Сk����k.�� ��~�{Qs����
���m�}�Q
.,��A#X���i�.���>ޢ�[�0���ٛ���g��?���<}�6l½ݺ�p^�e�6������X�5�w9Q��B�B�~p�΅(�B�9�d��L�௜�c+r[?��nC�����r\_! �M�/���1l�=����j���G`���Q
��
�6�:�l;�r�>W��'H,�XZP\O��Y������o���g�g>������b-��ي7�]~���E��/�>qI�%��W�X�]��0����#8@O^mu����[�[[�.�U��X�ِ�\^;��?�E�r�����Dܐ�΂L�LRg�(Vy�G�<����n�Ti���X+�e9%�˚�X��:f
W��l��aw���UG�,�ʥ/r�]v?R�4I>�f����8)P�m#tEO��fWK]�M_f��U`�{��pw 0��$R�b� .�d]7)0��"��Ͼ9����6��R�o7ͷ{��d�ښ��p庑��p46�h�����n�����1�>�߉+u>�%n��)U�|Zǟ<� (p����\�̉���KL�I+�r��j"��1�j��>z�P9:66��Y��"y�.2���O0�x/g�>��{�7[o��aTQQ����j�\�U���sk���Xp�֓+ ��_��7 ��E� .S��[	Wpl�h�`�0�Z4�.�d�;rͱ@'�%R����6�Z���@B_�]e����`h�zWr�~4��?�j�}�2�r��m�c�^��Ջ���D����=��Yp @y_Y�S������2��|e�g� H1���S��tЗ��v��ˮ�;t�d�P�!ϋ��M&�`���@Gg+a"ۓ�s~�}}}�Y�9 _o��DJܲ��g�z=k���+���N Dp�)H===�dJn�^U�N��$<�,O�8TUq�W.`kdy�# x����h�KrON='��<��^zt�?�D� �ĕ̫I͇��HY�Q�52�ѪBXOc~���TZ50\	{|Я���U�H���߂g���*NnJTǀ#^�!O��P�����,4�:�[ȧ����ewPϼz���1C�N�dHژ�Q�TF��'�ޡub�����i�����i��7��V;0l�f�>�WdQbw�tZ�>�s��D,S4~��QFZ^ 3����v�KՔ�=��%�L>cY��J4c����� ��|w��Hޘ$�sO�ѹ'*�i�[� �א�'x�1�Ve�ܤ%�P�h��ї�U��k���Dx0V�g�<�t-�u��� R�L܉�G��]ɕt&�GwgjT{�����QI!��IP��bƞ�:她�
�����k]�9�R�0<��ev"��gW�bWTn�,�s���G�#��q��ť���Y��55Ғ�����*�Z�f�
!s�X���	_q������'5g~ρ����r�8� ��y=q�@�#�'E� |:����M��[E��������\�{����������j1���pWh��X/�bo�uk�;݀�G���dc�CxLzn ~�R�,�F3�Z ��@B�z�!����疗8�L��f%qA�(�����NY,��)�k����H�}Y��#���ޒ�S�+}�]�N)��/�H2�K�(�6aͭ���]e>�u�ީ��}d	�B�a��R��y@.������1݃����<�6�L4	VR<��C1����uL5-�n�G6��r
R�����5���*v�b��?	���X�%4���yuJ�~�����?tt@�!�����]3W��ψB=��}r��Q�P��M�������5�{� �j!�d��2�RN�
⨩TU��?�<�h�V����2-��9`z(�Q(�p�>�l�u��m��T�W��/����L��
r�����qqq��@�ĸ�A���Alv��?.S�1k�ʃ�h��în����{��j:�Ӎb�&�Z�`ɜ&��BRŐ���[^ΆB�rKJN�thA�Si��Y�JI�"�k��t����QN;	���#�نj.���{���V��y��BFJ�Oʲޟ���z��!vŀ��d}{8Mz�pt,��'r%�x�X3�}z"e%����ܢ"F�Ǒ�`�kx�P��TZ�
��J����'6�(JQn�Z��_dp���ͪ��Js����sۗ�)���NKK��? E�N�{{'�v�<X6�u�B�I4 ��=zt����fVV<�e��`5�p�<����OXخ�{�`�L����X0��q������ɓb#��󛼋�T��M� ���G�#Wh�o���G)�o�T̿�~|��Cvv]}�" ��{Er�ͩ& ��M4�A~���NEje����!Y��z��Nq��m�6gs2�1Y��2�5�0<l��V����th�K�e'+׋9C]�o �{5r	|^��lY|)(�x�q�}���npddv���G7l�Y 1�Ɵ��$�gѾ���=�Dl�M�21�{�����5�4��P`@��KJ�}��T�X�AQG�K�rS@���UZ�A�N�RB{��/�1� *25�,�դ��g:��{{ �6z(Β��w���]�0�*�?q�n��!63BeX
5q���{(i������<k����;e�Çۯfgg� ���+��F��>F�9����XéW�W��B�>�l���͎D+��L���̫8�?Ըk�R�F��wvv���)���Ѯ�.e�����;22�A|��=p���99j�gs�,٘�8�z��ei��
1��(�C3�*�;�
�Ѹ*8�+�{mW�`����d�-,8���=�x2�TŘ뺰ܚ|���4�؅��wB�߻�`�Õ�v�H_7�W��I�&^�.KHh��y=�LL��Y�2^�R��2@��"c��s�mAJ�������(�l�o�C�E��G8H�"Yd��i��_��|K���j�d��
�b��;]a]�;vi:��D
��� �&d�>�S�����`<:������*++20(�*�Ak�����_ĠذS�	A����N/�Q�{m~ǭ�'�j���8����/��-�� �fr�*��M?�T�$tg�p⽸�_1E�ˉ�����BܦX�F��9���#�b�~�i��E8�k"-0��񸷡'��y��L��z��>#1-\�D������.�FZ��˸_T���6` ��"LL6� ������}�V�;��B�\��~�: �-���5�Jz��FzPiw���d��:���8a�QX:֓� [��]p���N�5O��p�z��F�u[6��d�n7�53kSBeY��6\\�zs7�d�=�,V�J�̊c�ā۳��Ml�$7P����T�<Ԛ�,?�U���W@�O���@����`�
'?^�V�V!��Fq����0L�$�f$z��5}�>��ı
b��g����~��Z�9T��c���^2����\��ؘ�r���
a$3C��re���0� ��fR"�72��d��`��Y
�?�����;�M��e!�@UHDU�9ٕD��R'��m��z��+\��;�BAG�v�����.R�>U��h1�H��P9/nbP���Q����˦���a�#xz���h��	�L��	x|iP�zP?m�⦞�͖��f�I*J����?O���j�9��Ob�;X}X�	�y,^�yWϿ��n(�n���99X�PD�G}-_ �믖ӧi��6�y͛g�a@V1�f(�)P+?[�K�ʥOkõ(�V�񰌹���	����b��z���"��x�8}�ϲ�M`��6pKD�`�qNF���A_{
�d<�K�/gz�.��� ��ʐ����yr�Av;=�1����e-�QiƢ��X5�4L��.+����Jt��U���׽hĔ@���׊1��#�:e!�Ӝ�H��8��՛���1lڻ}sAu#��B;\/�}�C��k�S��J-A��Nx�e~,��[��zL�z��0�Eݰ�<AxNW�7,������d��1��bN 01R^�a� V����Σ:R� A���
�;�G�S6	����8��üi�'z�G��/��Ќ��o�R�Je�!�;�� s�� w6#��cb��9âV��4�����)fL&B��2OP4�a2��~v��Zqc�<�i��$��B8ON{�;8_����333�:Z-1�O����_7"�3��i7˃�x���{��B__���!���d�O��جd��s��T�H3#�ܔ��K����aNG������z��7 ���i���H���o�-3?��x1���n��$!�
ӫ��,��g�v$�՛�󪄳��W���Gg�/Z	콧��������=!��{����<��,��ȴ���=�V��2Z~c+_i�*��XlP0ڽ�����㚓~�A���3�.gі��-<*>�v�k��>#]E�n_Іĵ �%Y�Aa� �h5�2���qA�0�V�m�׮�ax/���Ӽ��wr�~�]��,guP������G��"�s���ey���Pʢ�a�5��q�~5����M�ʳ�aJ�:q�y�\��	�sj��}s���8����TE��m1t˞�1RT�Jk��_th�27�pt��3Vf?"���VjTb��;�=WW����U�ע6��>��`��:Ҡ�7|A�u�� ��J�3ˁD��D߭/��bCL�/4�����<�SRx��B��m���[=��O)�O�&)��oWx�64�^��`�ts��)�m�u�4gN��R��IU¨�>ǳdW?2u}��� ���"..T9h�LƜ�@��I��!�[x�)�IS���{�v�mj�n�It�Q�-� �?V��q�)��}��TB��~9nu�$�9u� oG_(l4#�|�� �T���e:�q1��۞v^���f�������Ey׉�����Y}�$8C.K���X&V%�X��C��� P[�ܛ��}$��<e>�w�	��#/�jHe��'�� ��#�)�)2�6�#y)��C=���"���F��=1�7H���|���r�-�Uk�{����9j[�r���G��A�J���g	B����{ƈo�j(��RT�<��g��T������ UJ��*A�#�M�OxСy�/��\5C�%0������b=hmܾU!��P�Y�e83#1 �U�<3�FN����$[}�a�pZ�q ��CX_l�:� �0��C֒���,LW�R;yU|f�a�T)W1O�nN�&��.� j?B�r�b9}d�G`��k�s&d�{�W��	�<��C�'g�X��nD���F�s훟ٽ{C�=VI�VI^���˙��GyFJ&�k����g�,��:�5����d�o�$d��d5�Ŀ�s\�`XI4�/򺗧�0�����0P�����������ko�b��Zd��eW�o�.
���qA��N���>�����a��P:p�������Z�8�H���u����\Nr�� ��ۋO��<Ɣ1;;�.g�7n�����Ü����Բ�:Z���v:Gպ�����&&5�}Elr�2�]>�����G+՜�� 9x/J��)�h䱟 �y����>�	� K���.|>��r�\�E��r�>}Ɓ'XØcEޕ:���VV��Vр�i���¶ɐ�gZ�L0Ԝ������j,�~r�Cn-(<�������r�666�"XxC���p�)%U�% ��!ItX�u��Z1Z`��q�8%6���l��hӈ��>m?����_��ɀO�O���vj��1v-�d[��L+\+ܥ��1VG<�������'=�*�U�7�	�n�R%�^ �I�0��pu3����f1�^�PY�0�O�*"ȋw�D6Tǩ�l������j����M�Ζ?rOD�W��u�Wx_�1澿��:�y�+��==�\}��yY��'	���}?��p��r�Nd���W��9処M���u����G��W���ǝ�7���cD���Q���k�M�'�̎���ΓQ��4�ZY81�B����o��A��(W�=��B�I����`X,���;9?�n���X�<�7� ����]-X�q)�{)�4��Չ$Ι�u���o߮�o�V�Ux��IZNO�g��G��ߍA!��f������cU�v�[)�vT���mi�\�&����:v$���Dx��7Go�u`Eq8��K��G�^��>?j�U:�R���Y�71Ev���B�����N�͕L��s��%F���U=-3�.���r����frPv���G�Ծ��ur~1��K`y~@n
�Փ����-����y�/�(��qb�R��Zf�T�*�i&#B8�8�V��K��ᭋ�%tt�w]�#���kĂ�T�9�wS������s������ťa��m�����|�B������Q��%"K�+�i�ܦ��@sȒ8��ߩ��ZK� af?*�s캋</%�e���%ғ/�x�f��ѵ
�7P�D]�Y]��i~�3C-�����U:��$o��Ͽ�p����L���?״�W Z�f�f�IP����V�h�[�*�1M�*�/�;�v+=�s������- �[�#����;����9�9���E���Y:�Y޴j����E�]q:G�P
�UPa���L�vPm�wl�	w������XSS�ObfcS-�6�U}�+kY��)��Aa�)�����p1+�JAEjmC=�hH��������p#[G�\	�ܿ2<+�U�F(�qS1F�� p|�{~���Cs�?�U�X}��m!օ�lLN>PUUM�8 ��ݰ0b��w����AA����vl�o3a如�:�����Y��?5#�<���C}� �B��������t9���%��+h�>��'�z�*"�(������1 � ��`�����7�Р�)�|�iJ W����,�\T�j:Uhp�Ճk|�H���Ĉ?��j@_�O �m6J��Uu�/�v��w:Y��h�.�(ׇk�I����|�U�� ��M� �+��h��fܧ&J	�*U�j���ϥ���Tw�l�G*� �<� ����o��\���I�\��u��0B���c+#�a��|D:��#q�`��'���*��v�t!S'����>�1��D���h���sP٠4�
��oObm}wN���/Z�Ui��q���}������(��hĲ���SZ���/�:����^}����{��9�4z�	Y~������V�a���:ԦH�>9U�$�10�T� �ˋ�i��v��}�AY�q����sgϞ>;�t�߬�S��Ā��-0�o��&��^x`x��3@�e=u$sM���ʎ�zw�~ʚ�'��Y�3����7�H�.;A������0S��4���<����zxQK�+�����`� [�98פ���P9���#���o��������R��W���
��ԉE�Z�������+����%qn'R����Q�����m/k�XWt�w��zp=���;>��\_�|C�6tƈ�;�XDM��ng��u�i��i:�h��/�쿝�qr���ƞ�d���W�j|�A��2({�bص�����;�x��ʉy�NLd�x&= Xu�������3P9�x�����i �RR�ť���q�(��=������q��s�v�1A�K����M�f��)��I�8�}���q_�"����Ix�l�`�e�5>r9���*m��5�.?�G�b�{���K����r�,��-�{�o��PP" �Bus�x�4}N�û��'S,����j�_� ��\������o�w��9d�t�ϟ܇�D����K�	�I�zS����]�N�(�s�j�6�fٛ6���,xz4)�+�r�ޡ��X�V��?��~�=��[��f_�L�^�y��q��0��}��. 5\���Еw��5O�(e"��]:
\����ڡ���B��cl���唪C��o��%���~u/=�l���A06��!�u!�[�����s�m�x����}Q���l!˵nT�¯������;�I10ͯ����?F�0�1T���1MP6�Ia\�{�!� ����X�+���������ɀ$����<|��Tю�UO%���( 8WLW��*Z�/;<GG��^X����{/w�]CM� x��6Un����96�;�\ɶ��_���_��qqA��p}�]lo�s?m����!c8@��7�#��a�F�.
1�6�t��*�^]�J�zϟ�8�L6:L���e:77�]��ƶ���]���J_�F��rq%���9_ƅ崋����c!���P��R���h+�	���Z�VW�]���l�d�6	��;>�n��}b�EcTZ�D�y �W���ITls�5���{�
���̋���N��0�%���0g��#c҅&�]����r�U�y��Y�>��l�b��P���3�|,���E���̭'�����zI[�� XI(����O��\�l���`tu� [���Nk��Lxec`k�����Dj�Ƅl�^k8�*b�ꄦ�qUQb֟ ��.'o�iw�dw>�"�4
��8{�7�c��)��4pF1���Ba�����dՖ�Z�;���DV��{��Z-�DH烳�o\/����d
�p���*[�֭d9�(�yl�5�ʵ�'�	���2~�2lj�N%��T����/淬�2��X��/<#SI�Ҋo�xw������?^Y#�G�!�G�}}��CU�ӧo�ۂ�9�̚h׆�{w�?�.Á�u����։lQ�����\<����g�p�(V�c�8q�I�IZY^^�}٭�%$�װ�88'ⵍ��H)J��e���j���t��RlIdǠ��f�[T��ļ�r���c�S��h���T�nN��]��yf1���u���ɩ�w�!p��2�^nnn��! !� ����9����Sv�����A�q��$=W����˳���]��#��s��q�5�\S���u�"�����??1>���l}&�4ޚ��|�t�H�I�
�Unm�3��#s�s�P"����if2x����2�w��r *M宾d�iA��
�=�k�Ξ�d��DYƌ$�s�/�F)0f����=l%Gևs_ ^#����|6��MM��3W��3R�j��~� ��Vy��0��^�5z��~;������M�l�\f��Q�%��t�i�uN?�s!2�ɸ��κ�-�C�ǠCD�$�n�KD������%��ߚ0��x���|	@[w}۲�k��6ZN��̳tCq2� ��%��G.v�On��E�����J���xQ�4 �v���u���e{�o:yם���*�l����W����Q���W �"�����I��R2��.|\__?d'�G~�bVG�t�-�,^�(��(�����imA#�H�m���ha�G[�����}�QK9�N�|�r[�9xEK���"����ŷx|�SΊ�����!�n?�#�;�[~� 80���Fhkiz���S��piy9=�+S+cX}kI}�)-�[!�����C`r$v�b���əO5#��H�/�y|��N{b]#�W��&��!��,��#6sy[�XYeO��d$k��&���U�S�ڥry�22l~��!��A�h��[暖�rX������hX0�h� ��9��It�X���O*���O�b@(zh�H�i���{�7WrjmXe-迾e� dJ�ζʸK��W���R���숒ܚLz�?�[>�'!ܙc��Ԗ���gf9G�����!D�x���G�T�8R�i����bM�p��N���� ($�b�Y��C�˾�)���f+�b�U��>O���5������n�}3������~���ۚ����!NW�/-Unvm�(��Ŷ�g�b0�Z�O���g�'�Ϸ�:�M��2\M�c]�Y���>u��ߌ��݃�̬2tg#�&+%K'.�y��y��i��ѣǎշ�(�����Us?�Yև��>+C~#մ���_��7���&��J�?9�ʑ�L%�S�����z�H��U�3O7p��D��� �S�f��~���~2�b��p$%k�BC��l ��|�7���%��s�x�@A�ה����ro�}��9����''��+
���{��^�W[[��(��jåH��$�|�n�=%KV����j�8Cb��t�y���)��`�1��@��u{�����=|r��sn��E4�~-V�7W'���������2��m�c��8%EEM����+ws��+Y|��8 =�ϙIq+*����no}���NirV/�X����j���Ԯ��|��B���3Q 5559�}���M}O�����x���?�<_)�@TQ�m�Z%d�m�z �x#Î.>�Ǘ�tXÁ�$�������S+o�=��'1�٠�I̲���h��s�K�x��k�wQ*ɒn���S�P��7����-�$�g�JC��Y��`����/M�p$�	��U��M鱅��fv����V��D���u&�ω����
O}��[�6�?4G'*phn��x���۪��R�32x:����G�g����y��Ճ���n��~!{hD2إ.�m�o!���6?���B�U���B3���Z�^�OڽG48k ��`����I�L�}z����J7v�:$�K��,p�aMb�������
���u��������+�)���#<ޒĩ%蟦]������?)~oD͓�����@�w&�ɖ������a�9�Y��� `����2=0������9o��@n���e ���tV�@��B��G�Z�_���[B�^l}����x�9yf�0��q��%����0riU�u��|D�W،�C*�}��˧Ad������#��v���v�#�|c��{�K��Q����V,��/w�;�E�{�wVG�e~,���I{�@ �7F]hHBF�o�@�G��I��<h�L��`ao��+����	��+�>g2�AFhS}��&���d�����K�GJ�v������%�V�L�j;|�l(�Ž;����\���V���q)�@zU� ��޵�=[��{�G�L���[�L1sp�x_f��$w*Mf��/��^��(�9�H�w�Y�(-e��Gr_O�ʍ���Qc0�������;�omVS�_�*)oS�6-���ߥ�Ǉ���Z�r���@�3pG�ưY\R2�-��3����A8�˽�tL'S۬��]�L텐�#��_�:U�Q�\���CIDbڿ��<��q�jˇF~0-�(��/2H���u22�n��L���d�C�s4
���f#�����M��h?�jзW |��aY�Z����G-��� �?tA"'�ϊi񡣕��[����/��`5�h�j�u�b�|���th���&J�(��xz�A�芊���5��7�1{;f����-Ҋ���T��|�nWl�+ǡ�CsM���T��wW�l���z�Y0�����#x�|3�d�H����y�Y���R�ou�sǝ�1�9<��S�<y�����Y��z�z�"� ���a�s ��4M�w_@��<M��wC-�V��8m�W�V�Q��e.�r�t��9p��a���� [)FBpW�S	���H��e�x_�l�H��� n�)VLTR���3���ڝ������AI"]`��8���/4p��<i"�u�t�袍�n~0�H�d\��{�nkG�)�����	�Ť-�Rǝ��m!�?9}r��s�����"e�%���v�ن��@���̏���&;)��e�3ʀ��S+v�X��"ZP��Hs��Ү��6^�����LTB��0�K���.mPm(By;�n��^�}���|����J5V�qz�R��#�t9��B@�])�Ǌ5k&���;+�L䑂�:�#:�� ��̌+M�?�^t�PD�ɟ�-�+�-Ҷ�{G�Q�8�C_�����\ q��X���5�]ށ̎^�3��c~�v>�����}.��aҾ��@ߔx��SBI]�C.6o޽�����`Y*�*
c��M�����ܟ4��bJ�Z�0'Nw��y�e?iF�?�gp����[�Ϩs	�V�r|�/�������埡��ZTS����W�����>�h�;�=4yD�f%��k�hΫ����
���k8���o�M����ghW�\"��fg�U�����!B0�;Ƈ�%��Q���ސS{T��/��$$�% �qx\�WX����j����H�F�O�tw��B�m��Wc�_���x~Ha�D��U�|ct�`��+Z3�v�|
��v	�T������C���U�~�  �
A1[P(<�����9Z�p��N+~��J�Oy!P��.ZxQc"\MW�� HFp��ŋpL~O��ℒ����ާ3LMG�18aٹ�d���\����3�_��s]}��t������Ӊ>����f���ƑϯΖX������;�}Q � a�G�*wC��Z D{��8�ҍ���[m���\'mm��%s����~���!�'��Tq�pPu�_~E�ޫ��7��7���&�r|b�ҪX���D �;�O0zL�oN��ιv{r�2"�9�6�����5g��+Q(��rXȥ�|�wu�5�18@O�Xv���k�_������j��d�s��U8 �.s���I�|{�����΁�	�ܽƥr@��V嶬�\w������-���H�p�ߙ��r�8[�7�E���3�7+qi���Q�E���z�=<J;�jgJ2�/�2Ρ�yZ�:��o��y��}�����G�.R��^��^�`���ʦJ$w�m�`�������i1�<<�V���v��~y'�����b�l\|G�wF�P�p�I�l�"��R��R�����t��*Z��߹/j�<��kb
��vZ���ӣ�"��|y���E��^S�K,�
��o0�l�n9D�zmw�#CK+	�LOZ?������Y�F�s33*|�.�����U��%3p@$n+2��u�*�G���5)�V;ݽ��ֵ�S8�.;_c����b�<� <�����@��@:���W:�oL�>�W#H���.^����� |W�p����� O�����U���{�TZ�@�.�v���N���mX�>R�h5{��CƓ �L-u���Op��w�v�W(>�E��=7��]����f9�y*�V���FǕ�CM�;�&24�<fŇ֒,�	=&`�;�(�����K��Y@� ���\���o�ݟ,Y:�u�LV���P�Ğ_���,,,�p�>&����7K0M�q��K��a��0:����~�	Vr���F�8��:��Ud�֣��� �!��ϋp�E�i�4biQ���S�pb����� ��?J��W��ݻ7׺�}S3j؟�Z��%]]ݥ�eE�/xtH�ukq�X�du��aq_N�qQQ:�H@E� Ą
�����7���P�r����b��b|v׌�ЖY�2<ɏ@x�R�T'���?���+�V���1A�[��V�D,ew��Ѻ�IX6����4�R��ɹ��lF L �������ͅjh�V�lUUUx
@@׼�B�/��1���c�ok[,%)d��Y����W���x�dr߶�/G�^�:���e�O�E���x9��A_y�/��E2������f_��C�K���Q��'!'�)dJ���U iL ������C3o�L�j��S�0��\�`��Y\7�7�q��-�L�mO��V,���7�s�J��L-��Xx�+��;�)�>-'\�󿬺�kS�3P�7F�Z4F��js�bs�B � ��V	@`�%ɲ����`C���*�P��Z���@���k4���E�̬�q������"t�N	��
�<�A�|�$��`$�0;<�vV�&[SG?�ZYm�˅�u�.��j9�c�����Dw��g�˗�$ :�?tb�d��(dU�7�N�n��l��)�'�W�4��6k���<X�����iW2>(����k�s�9�5�7������2J���I���$VU���$ao�\\L ��z��i>�>��jb�2,���Tn��c��k�pf&Dz.歼*���O�W�LN	�H���B��i��,���U�>��o�k���U�~����-���s�ӽ�À*�NkR���Mg-@ӑ������k�X���m�0�ui���a�Q�����I�'$�3qs�\��5��˯����?���+$��kVwE�X]�'�g}���ƨv�IhX/���M�>-l�\>Jr���	{���(�EQ 6 *��HxĬ�퇕z`P,�0�iT�W�A��C#����x�	 �BF�0 �X83���W�;�ɳ��"����2f�Ջ�e�3:"�Ц�~/ ��	BP%��ͤ�E�z�Q.��D�����@�u3�����֕�Y���pt#�%���L 4d�5�;��ǹ�!R����b"{�!j6�r���'����0L{�aS~	�=�p챈cyt���y�S��m1d�co����O���	�mE��~Pŏ�� ���1P�Z�C~�!�Xw�dJh������]v��=��D��D<܉��a�+U���u�dX;�"/�J�Q�F�ηR�S�� @'����˷����!}Mfe�# ��->���m�_�}���-����Ь�
)��y7���Q��:���u��g̀.�#G�i�.�ã��eb����� ��= >�'t>�<,�>S�+<:�4����AQ0�I+�����E@E�� ��?%���ĕ��͙��ϋ�wtǤ0�9TA7\��� 'r�X6���e�f�kq�?����ˑ��o�L�i~�S��<4�"��b�F�3�	1��%m�&M�?��A3�*j�L��a��n�X�N�v��%�%m�/��1&���7��P�H�@N�LN��f�{���>��F�2A(��S�q��-������ ��J�0*�d�ޢ��g9�1��%��g��#�e���	p�!@��K|^�D�{}Exc���*�m$8��ݖ�V3��������?S18��	m9��8�[��(�С?~��D:	������"�Y��hq��G���U���� Ѝ6�++�O�Ő�q���('Ė��|O�/9�V�YO����d�QsҬu��ǜ���se��f�I��I����o�9Jh��>���ᾴ'�����x:���6�+ײ*a��0��v������R
g�y��Q�s��u;%<�=Ie��,f �q��x��F���_a�k�?\�T�K�?�5@�DJA@@JJ�F��<�(��!%�tI+ݍ4H�4HwIw�;�>��Z�Y�{�]�93��'�왯�l��<X�O��������0Ã*��E����s�>�0u��?R,����>�{�����t�2-���E�³�p�â`�%�p�,�w{K�E�xa���i��Q���6�^o�)*k��[������b�����z�������ռ�ypWO"*�r���M0�n�@_�:�͂�[$�B6<XY�����'�����w	�q������b��3@�0Ir����n>��v4�u�=�K*BBx�X?��,���~/��PVi;@�����mX5���[5�%���,�n�s#Ywt}���R�3ƾ�q�-w���+K�Ò�@\Z��UE�?�*��k��jU�����Bª���� /����N���;L�M��vl���w݃q����x�]I���֫c��a5���C����Os�I'.��Z~@�.���뛪������Hĸ��K�d�	���9˿ҭO�r��i��.'�/EiOV�B):�+�{����%N~`�{8Gyi���2�<
;"��{�@������i3�-�	T��ۏ�r��?��[".����V��պ�<���N�\�}���D]=lTv���}��uDgə�,ܥ��?n� �y���/���b�������$<n�M�^��3���AB�M��@���"������u?���fY Z4�S+gp;�wg�ۍ,�����C�\��lrkI�8�o����k��o��=�������Nr�}ᑋ�^5[[�f`P���mlX��������g�@�u>�c�?:���9Z2
�.b�hV��@!���������_W=��@tٷ~)��#78��O�ة� 0C��:zC9ʭ���E%�Dtx�������߻���P�>�Q�����onn�M���.3VN_��\<V����R��l
p8.�:��u��Js�xg������6���I�!4��'�ƹ��fkm� �'��Mw�]i �&�?�N�0�l�}u���n�ߣ�x�Xg�o��]f��[�K��,$U��2~�#F��rШ�>�kB*��X}���(a��%^����)�I�s�i^B����_���P�kwF�;����)�����3[��3tV��v�97'�V+��؁O��Ҽ/�,rN>�TA�nT7&�q-��P3wA8l��w��J~���V���u�  [��v��9n^_��`��P�<0dt�HԀ �6�!�C����=K)�ҭ�����є����V�QK[���'�MA���ӖfL��<�����6��Pi1v���X��<[�2�Q?3����W�X������t}������kL�X�>�v�, tlZ>�W>a%N)Թhu��~Q0&��S¥�&w} ,F"���tmދ�|�s�@�Y�N��ݠPx�;�`��x����"�B������%uy�~�m���Y�D?/d�%;�)��Q(D��'�ͧ�:�?B����.x&U�*�[�b4ߞ
_���3�]�[7���]G�$č��/\�¹zFvSB���L=f&q�'��������P���+; n�3z*�.�H�6��Ȧ	��'}���2D��f�\��6U@�BI���y�3�����%Xt�ZM�m>s;�꨻A��I���t]y])�Gݹ�*��eV{�$?N��#o�9�IUW�C��nC�7�rs�a�i}�� �z7W��J������-�I܍�ʥœ���y5J|۰I8�E����N�Њ(H�~�{�XS�)�%�$dz�a%!k����2��jjN�ew�	��AjR����d��b��F�ۆ�>k#p��\;�C7݀�O��\��H~����Q�ʠ�[����p�`e�!�I���>�nB�e&od�~O�r~��&���ʛ�TB�3/Xo1i;�hwh"��0D@B@�g��T�<Z ���K�����l�6��H/��죮�B��F��C��^;N�x0Za��i�ַQ�	�`M���h�IOg+μ��y�F� ��k3!����2���-��)6 �a�ǃ s|���Xe=��@���pږ���X�@6vo�C)�S{���vvs�<��|g���應G5THHHV��l������*�~����:��:;;��� ���ic���֗���ו�d4]��DM��WTr�a��;l�Q�qlIUx��q�=��xS]-$-���AW��O0{��M�ʚ��ii���\����a'���b��ۢ �>k��fPV���V~��K���0�c��2�Vf����O@��;'��v=j��y+��b��}�g�#���� =9o�R�Ud��|�5RZ�xz�:9��Q��E쾋����:#�jP>~���6�=����`֣��"��_�x���J����S�-+xqq��.��4��܀�$�����=��������V=#��q���g%U��g�	Qۏ�S��%͖�y��ۀ��Z#r�^������/RRRv �����!�~#=P�����#:X�FTƟ��e�l�.�[�]/���� ��
���W�:�/���m�ԦsC�|�н�ZX�������J�(�Z��k^��g���������t���+`!)����f�C*??ً��.�q|�>�qT˿}����S򇯷qe'|�g>�R��e�2�M7{�<�?�X�)900�Ǚ�a8P�=<Gijz��.:��=������+��?=<�cb�I.%�e%.��%�8��Z���p�N���سw2�OfV�lMԨI6���i��3G�ʦ�@�d����g��N����A�~��T�|�Է�2\������c�._��%���ѣG�蟚o���s�����wQQ_PSJ����Sj��~ᴦ���ÑF�- p|�o�/�q�5@u�g����N=���޽K�X:���	����^+�ƸQ�\��Y�n�������~YYR��]]��v�����r�h�F�V���Ρ�]]�&V�����
�>��4�M$��HII����JYP�aN�#[�sc]�h�CB> B�622���q���E���&�fLL����ΊtT�����3v��߮m:�~}�����=pJ��3u:���95𝜜���|��t�ҭw���E_>�66A�����9K:��,��c��o-,`E��C�h�ݫ8��h"RR¢���\:���������e���획���9�=�� E�1=f���"�Y?h�*��< ��ܔ��;wHiiŇ��o�RW�G��>-M��ull�������C+�MF��-��؅��q$/�雁����+��C@�nr>Oru?q�,m�Ŭ��	==��43)ٮ���ވ���L�~�B��m�]
������W*��8rl\�7&''c�վ��ǯ++G�=Z�������8ՠǜ���Mz%�rrP����[TO��H�`���ݻ�DD�]1��(((U5��X���敼k�����z2x��������S�3�dj���^���	����P.��="���ݗ2VVŽ�����
����ӑ|1�޼ie���o���~�~钚��꘹f��{����=|ghI.�(  R�ߕ��((x''�	
��n
�{��j6p�5��%��c�R�>S�0F��e�E����~)�s����qO�������^��t���t¢	���OD��VX��ڥ;������n�����/��N���U�ժ�S�ⱐrǯ_QU�"��d��Fh�!;/c�#0�^�}��g����5!�͉;饥,��F����UԴ�M@K��F��l	$�٬�2�zui؟**"!5=4��m[s8\OK�8�Q���T|��Q�3P�ެ��o;"�bb���V��$#�{5<Y�%�qy��Wcc����I�x˛��_�z������2��+a�-C��HI_E"�c����n��B~�K�&༊Y��XR�o�\�$�1�����z�|h���$#/������f�F.��;r
�ssт�N3{]88 <n!+h9����E�Y{�w�1Q��>�R��"+++")����^�-��������&������O�݅vE[[ ;j�M�����ϲ�bd�TVVf��4�ݤU���9Y��pFP2�p�H'	���aV��5���SaC�
�c�WH�?*�$@��.�]^	Ivwt�ݖ�E����g���v��K�^�6~VS��Dk�����Z�/Fܵ�r8�ns)��g�g��K�VP���/*�
�ٽ������U[[� T��jFR���A���#m�5s;�F�''�.��i����u�Bh^3�h}� d��d�_K��j�ӧO�_�ĕrp�wg��p+ji6��#�'`Ƣz<%����N����)O�'m�KM�J��1-n�tt�|��\ �իW¸Zzz���]���C�����SR^G��H�sx C�-�wl2Z,��^Z��X��������0pD��Ӣ�ޚ?o�o�YY�R>Nq��6���ť8ha:I���������ْ����`����w�ȃ�&}�g�)4H��w���L��
��|t�9ź]��q0\+��
��k1��Qs��2�|y��]���䑑�t ��iwq1���B���@#ql�*�t�f��H��h&J�!��"���.0j���H.�o��@AEE�Ʀ��c�Z����G�PQy���Y�����o�����3�^BQU�',,�9@DÓ���G, >����v��n��5Q*E"����d���g�����O�j�3@�Y�x��~�u�WȧɓiN���;y������9k1S^A�w���[��a��l��H$d���2��uT�?�Z/u����R�r�����.�uzw��:��W2����x&a}v��Ǉ�rλ�f�D?��\�=���er��P{����?�ͧ �B��0�z@Hw�D;͍�	��2�S��Z6��̣�6h%(���&��6D��L��̜g�ؘ�OXx�n����Y	���e�j\-�A097��l�Ez<u�_�~�6�C��u�P�.V�V]R��^IN���e�0�CJ\�ׯD�U�̔>ꚓ}�&��zرY?���o�"gf�����orr����M���]���=�^ɣo߾�lm� ��%���1�U�mmw==N��#�tު�X�
�3+'<9����gA���� �Ϗ��êwv�W��˿:;����u���@aҭ<Ѥ����**~��"��n:�]u�ŷ�%��ۑ���N�%@ �,���D^B�ћf�|�yFD� �.��F_mjjtגW>�=;��|�q�Hʴi����XjBF�PpHH�e=PP�F��^�Ө�]�6[p��*�7]�=��z���5w�8���1�g���#]���C�"���	͚j���mY!���"��+9����,=�@|��>��#Q��线"[���E������qWGH���|Q,-`S6,�e��X�5-��+���tt-�^ )݂�J`�;;/�-��+(������a����V�䥣|u=P����D�z���4ᴖ�����11���}E*��p�>�1���677g��
�ۗ�R��3��G�yrv��>6,�v����-���yjT�6�Zpp�?F3<1Z7q�p@SՒ}��){�����Z�O�PU`_��Pj�X}0	�9,�N�����h
�����9.h�� ����{�n'a�.S�},�o�X��l����spd��o^��!""ʓ�H��/H_���3��l惎N�4;�&f'��	@�>�2{��++Y���f���.���{�~6a�^Nr'&q;&��gcgw�h͍u����k]�&�9Mwm�˴��b�8XDӢ��顤���ـA-ӝQ��Q���������9�=X�נ�g���V����+�JL�a��}����%���������=������LLɆ���G ���o��s�𲭭m��e��<�e���	nn+����u/u����$�*f�т_��Ztb�ۯ.��i��z����N���`��)=+��	��aIR�Q�ѥ�����!c�CB��+<Кg(��ۛ��TP�ThA�n�g�ffe�t�PԱ�y��#�$$�'{��#̣�Tk�XY�����*r,��C����������/�����P�V�"�7E���̡�!q��k8�igϴ���B�eӖAE����RS��&X��wW"��������G~��l"�9��EF�,����F���W[���OY̩N�'�E����+�Uݹ�TU���������%����:+��/��!��F�ꬩ
x����&+�8�[ﵢ"�R�ʷ���濾�i:k1+?��*eTT2GO���_'�7�\���xz,%��\A�K���Zi�y����TXw��*·f�������ARβ���󋰰݄��'��O�C�#�yh��i��n���v-�v-?B�~���%�<�#�s�2�9��4��?� X+���y�{e��+!g1�hU�����P��}B����y�d����Pr!�1�냉6&e�4�
_`V��q�oM�Ʋ}���	??��I�2KgE������,���B��k4�6����),�,$<����~�\�q�U4J����d��l�6��`b_�IwRNv��&7x�ګ���៵��J�ws�m(Wbe|'?�	&"]
~�P��f/�Vd�h������ޘA�ݿ�3t�|�����W|��*=IIt��)b�Y�,��o,��5�{�=�H��L9�1���E��}�LA��^ܫ���/�"���r&&�6��F�(\���h�)ng��+(eq�+,�����[�����H����H���e���7p~�la��v����}jN��N�=U����v�W������|e�N/��G���IO��C��3�(��h����������5Iq�X��ר�v!�$��#V�|rv�>c K�B�T��� H���~��0?/�h`$2"�	9��t�on���ƾ�[�dQ�.P�@ ����p�q�]��������6��U�_�Ar�<m�A �T�>6������`�·�[�������;\��-a�F	���3�0�//.��������* �£N��;��ÄN)�~� K~����4���YZi��H3VV`ҥ~�����3�欬,��ٜ�|X�~��뗞������ޞn�����E�m��V�m�3i�c��i�P�Ӏ���I�;����	?V�%��|��J��wb���w��J$=77}5N��	&&�:Ъ�$�HK�����il�vab���E��~"�bT�w�4�+Z9T�MA��L�FN�j�v �o@������iT)��+�6���5o|C�ѱ��?`��.�ɴ���no[��E�p�]7l�\��f�w@TTTR�k|�,B&�Ac��VAFE��_hb�ϣ��Yk����jq���r�o��8��yͻ<d�ˈ��1�����2���;de���4TǱ�����D���]���n�GDD(������pĐ�zh����TvK�ϒ#Z�U�8u��oۡ4���vʭQ�d>[�<r*
33u�h���X8�����ZZ�`$�E�����G�)m�g����� ��e�q���&�ҾS��[�OP�����iqQQ�0y5���^'���z����p�Y+n�����R?l0x(�H8Q����s�x����
��,,R�{�������|�N��FUDm� ��.7O��1 ����n���]��'E�&���2M�>�**R�D/��:����Q���j�^�����������nt������!):��������.��u�j����De���;7C�7A
5����i�m�П&��d�gKqt�[{�RI|y\L��	\w ��kW��XYY�D�|���!#�=�?jFF鱞����-� <~LSU���^��V@	u��q��,F=x���%���5иJXV�-a<�8"2�$If��mHG���/�M���G2D�f-�/X��ڇ͆���)m
O�MB��=�Z2�YͼV� ���W�i��:�f_�2d.pi��O*�ճ����*��j�-aa�!<a=v)_��D�?*�1���E�l
Vʈ�ʆ�	��f�-9#	��VII�0橔b�@��m�$~�� �2�I���1���!���%��2����/��V<��ͬf$Ei ��<=X����r4�a�V��^�T�3���&���.�# 򆣂u?�w�02b�[�t�<��ɷnNL��U �tt���ڊv9�����M��!=�4*�79��w�`ջsѳ]������;QAІ�R_��ƭ�§�&/5-�]���<5U�YL���2����[f�t��")}~$�3�_����ZL����X�������<��qpp��l���@@۫c���n��aT \�P�7]N�{H�j42����T^-����d��!C�$��o�J��<���S4�`��s�<G$��7=��~+�����2BBC��i3ı�����L�]����"<46�ނtDkYE�8i�FH�d�^��L;1_���}���Q������Lo�ǋ�r��Q|��z�`��)q�O��P�2���k��¿���i��N�T��r�K�'HJ�2�x���0�o[R���w;�yq�n~<uT�K����4~���$���?��;����G�x�({t��Ü� �{Xx8y��/�R��I�2"L��\�A��+C�F��	"���ïm���bd�Un)�N�Y<��oe���C��|��I1s��t��S�6-�xc�8]�P�(:Uύ���Q�������>qA��	�]�Ȝ�+z��^�
��b������ǜ N��}�Xk��o�p*�/`[GF������#�$�UL����u0�[#c<~il���u�tR�m�+�c�&���5L�}N]g��ß�Zރ<�+�]�>��f�STV�pt=;lX�!��P�	�g '�e^wB\���*t�����IT�2 	r>>b�iW�x)*X�Ȑ��a�p=evnւcƆ����~�����&3�!�c$4x�`?�t(���@������U�HdRR�'��&j^�	��KiMM���->>jҤF�*���KJ�ÿnM��%5��N���=8A(,�ݹ���	>��br>
6%5��$g;(�?�HFC#*�-'.�j�7g9PP�:�fWU����j�		�.��������C��.CFשÄ�IF�q�}���·�r��`�hi�m%c�'Fg�j���{~4�ht�'������-���j�A����X;�8!���Yҫ�~c/g�9V@N64��0X4�+�gѳ�*�H���}h05�qCUU���͍��,��Jv�lp�g��6�> Ŏխ[�����J�{f-���<�~Q�^�	0�^�1:���+���T]��Y(k�'CT�s�kNĹ{��Y-gbAU����00�������wZ�=޾J2$76�`h8;'絴t�v2>=����ײ2Ł���ĵy�b��da�z%���|}:��_��b���?6D���$VV��0����q���<"*).�����cxq�n����O���¢��JF�(���a�;<X���Gx9�	J��B͸��A�Υ�ԥ�F<^�޶�uc�p^�����}3N���HLD�%�ZK�MMM@(��3���kəv猖b��nk���3���v(���s;��(�aeЗ4�rq!�5AT6�/k��"���a{8�������*ۜR�#f�__���A�ڮ)͎
�`���k��|���j��S=i���(�N�	֟���895����`w��� �k� �C𒫁��S��xRA7�4f���e.9y"6$b<a�����Ɩ3s��;��Va4�F�M�S%��ۓ�]��3���uL3���4%���wܐ�8�c?�%&拥�����"�@�����蠙��+RRx���K�qi�#��_KJ��*mcJ��@Aӌ":����+R�m�0X��E[yVʊ��OϢ����'��!g�g��)�vCu ,@v�s%ܨn��]�k7���hݎ��y1Ry��l���=�͝��+���p��r��������\�����!��2����U���eQ_��-	��RV��\YMMM�����Kh�i�J��DG1�8NRPP��zzzj7!�V">G[u ����N�}
i1� ��H�ڗ-����oq�����999��幹ᶌ���s���<�����돦�1�;{�x���b�����ksa�
�����O�K�;'m$�ʞ��R �N[�
�M_Pq]��V�I�D�Z]}���ab����(1;;���	���IS@c3���tx���O��U[�3�4�-�Z3��U���!G���Z\��1>>>jLn�ͪ�ϖ��N�Q6O[�����,ZͲן�����F��yOt=TE��4N���ul�U��C|'>Q�"2\+��#$!	��^_]@D��p�-�V�@���؝�I�&Rffy��(���II[�I^v�4���ayw>5{����8A�wӏ�y�>A� ���>����hm�'O���-�����߿���fP|،�t��l"��h?JA~�v�kkk׹r#�����gf�h����\��=|�+LUK��>Kg}�B{x�"���(��|.*bvJJQ���-��FM�E���.p`��::v�<��m@s͟�t� �(�N�M%u�Ҏ��}|@Grv���&�P�[n�cSe�%��u{��e��߹��KY�2#��?Y� �%5�)����ml>�̵@B�F�v�d���-H�d�}CC>@c��!;�++��[S���L������ͪ7�hF/�PQ�۬�]�a�_��jj[��Mw{{(�%��ﲻy�����	)�d���-�.	����i�6�/��	�B�wGP6�)%d��4s��T��K~�4u~x��o�P�3-&2�f���䛓� ����"q��K�d�����n�b���|�\�����AMM
�u�i��||��PFZF�7ZZI�!!�s�ʥ�ǀ��b���B�C[��&J�8	J�߅�u+�K�2Dv�<�[/�]�� ���^�N�:C׋~mI�;%�ë$#[���caO�������#��y P�f���I3|;��.Cէ@�t��@�Z�`W�3�K�R������-����������m�,*<�Q�������.��mljJz�����G���$!���
JJ r���f�Z-��� Ү��K�z��m�4@hX�w�)]9��R�==�QEEE��%-��t��Z�%GC��O$��;��������h�����ʨ� ���JLF�߼Am's�����IG
����O#*c�_��$��/����Zt-,�;m6w2��g�YhE5ВMM�޿O)=���������t+���'w
`���F�wE*�R&�:;ã6�c1D��H����O̡������9^GQ���;,�E�R��!ѥ�<\��H?�/���l�J,#r�诣m���n�ߊ���U!�UU\��`���dX�u#��.4�O�΀�����J�m�����^�x�? | eunN��`�F�����e��[�<��*++�L��f�0S�Z[[��Oq��M|��$���I���l���ǻ���ù�TT�D��u�8;o?��\������nR �0��IRG��Ё�o�F�l�}T���$ʍުW�B��
kmmM~�Iu�É��z>P �з昗�"V3&\5�C��F����� ���<|��g�뙷D��K�[W��f�j{t���؍v�Z�^�H|����|�����P{? ��\�//�#��{�n, ޷O���{�����p]&p?���g�W�|����"�ۤ0߆ � ;�к܍�Z{n����6充��;s͍�#Z�#����s�wt�E%DG/�'��)�nV�c�}͐����	?��N� �@�mydh��G*g(@�J@�� "�o}Z�N~~��Cȗ�6��T�w��*�B��q�s���;� �&��5qX�����)��99��޿�V�#�ʒSR�	s��98`�Q,�]A�y׵�r�g�w���f}�u`]Yq<b���7Β��@Oy������x�h���u:�*:�tz 5 rz���&��ya�����p�M��a���3�o[�\N�_�:::���m�;:꿹iVZ<O��6�%'9��]��������Ԍr~~-�|9�	�[x�װ)�ǧ������/��6�$cv�������-�$l��>g���ǉzE*�nN.���֑�|�U����c.`:�#��?�:=�ZF>o�TV8ѝ�a�57��&&��R�W"J���!�F�Ɩ���<�{���	&v��]Łί�%��?/L�����J(�&�'!��(A)��f�ⓦ1����%ť3���}pwƎ&)�ϕ+]:ɭ�@�a歎�m`�,�'-8�]�!��ռ`b�<?w��l%j,/������c� [S�"�� d���r�,ⷤ��.�����n���&ͨ�u��f�v��@�V"��:#q���Ru����#�,F �� �
VN�Y���^$l����Z!����2+�m[���X{�DE_��<���g����F���t��O��?	NAռ6v
�4Q�~OT�J`a�s�)o�0
vv|�x>�I������[ ��V9����sul^FU�>G�@w���A����A��f��Q��;_���z5����T�#��qa��S���Bm�R�k	�W��B� ��dW�����*O��v�Q<J��Bӊ�������~��k�P����fbb��9A���HV��ӣ?������X�w�ӆD����}�b��j�q�r~m�|44"�%��Dۉ�qi������ȹ(�\���M�Q�yg��~��{<nC&}}�����q�*�􆘽Tr-zd�HM*G�G��a�o-�jfH����F$�)�G?����>���HGi����h%��^�m�훚bxJ����ZrS$�^��D��S���c��:�o��!/��ृ�ǯ&$<��¾�#z ] �u�qĀ�K]�`1f��o�JQ0��4@�'�_j�V �pه�ɜ���'�w��VP/..4 c�%1�T�෺��qs�݁���	����X�7
��������G��4�/^�P)�����gB�~*Ě��$��+,�U6����5�0�i j�uO:��/�Z����vV7Z@𽂪*��:X�Q-v�/��7o�+'X�� � c�n�SQ��S�!���u�#���ˊa�9#,,��F���N6*P���
5E��_~ji/�D�ؠ6[.?���_�X/��7������&����k��z3(�1ف@/>3q�a�������!l �U�RG383��-N��K�.{����=�W<�ǭ�V��B1A�i����\\\��P�(/�R+�V�ǟ�۫�6rr޽��stx��'�W��l��RFF�	�Yz�YX�z�3�ֶLVH.V��>5�,͕c�Ȳ܈y�E]���	Z&��SL��?�����

!x�i�� �Sc����Fb?�J��M�kiY-��ˬ.`��{�@r�>pxX��S�Rx��s��S i�N+�.��T`Xŝ���`l^�x���.?[[Q{�h�۟�Vٙ�嗚���V�!���^v"p����[�Z
�;t%p+;l�<
6���E������ׂ5&#�
kO���3�����;��d����I���������(622�^P74�
�L�}Nh��޽~��t��u��~���t7��/[.lH0p1a�+�.�^g����F��թ���/?��=P$Ä��-m���X��ئJjj�&&91;i��R~�2G⬌�+��㩢�����M���B�+7�/$��D��(m��r��NN2��00�3Z>�t7� ��@cr0�K6���@�EA	�X�9{���.FzzI%`ss�Ro�=���q:Y�ہ�:[��ĺ.�>'�KO�x�BP�����1!!��7���ad}ۦa���p���n���9>�(3??	X6�����<��gS��Z�Ĵ��?�(�ml�9e�vvwG��ą�z�O9�Gw?e����ۻ���	`��F��T����[ɀ��i������QpQІn���~��9����V���ur��`���e �=��9eX �U6ﰰ��Ԏ&vOϳ�/ɒ���<����#9+KTd��������Sz�g�#��ã@����
J�s`����Q���&�Ʈ�F
}j�'<�B�j��qTH|8���v�]v�����5���ź��@�DHd���BxP �ڳ�>"?�GKn���������~��X��xx�r�S23E6@^�=�]�+�%Ƽw�^��q�Yy
hk�y؉	��i�H�1�2KKb�x�W�+��66�������4��w�?�����A&#���m�����
P^�k4?26�)���Mop�	���ί�W 1&PL@@��b,$*�_��Cl��ĔlE�����~�5+lt)�H���n{,�yb��<` P-`۴�Z����Ϗ�AQ �U��2��@C{��a�ld�'��L��fl���x/������uC8�쏐�S=��D�C«�啕���<D�r�6cY�mX5pn��#�n�~n�})$�aZ��!�������Ma!�Ģ��S��|o��q8l]gbi��/�`漣Ғ��'�O���3o��y@��Z���(X�q���HR]��R��^�4��^G�@V�bg��-�qMll�͞zh��iia�T���r^}�&&��<��Z�6�R�Teee尘�16>��[�Fpyqq�a�
�G�� K�W<ϑ�-X�]\3�-A��H�����69BV�_Ua��ׯ_��
��ePPR�#��ob ^Y.���Z�\=1��7P�!7�;::d���Ѻ�J��N�w�d/�?8�i�%���q����3k撘xV�5�W�`�^���3����4��H�~]��{���ťs�0���C�X��d3ɚ�Bm�K�KL�`��)X����3"b��W?�lc�����������num���_nЫ}i'�40���Q赆�<�`A�}A�I�!Iq���4����=�C��|*����A"[`^��zMV�Ӻ9���!y��+�[}~:<԰�0o[{���2E�a�Ȉ���=�������r�4P�^��s���)I9�	����,tq�C�D���N�[�����%�N6X��۴��3�|�;"imY������DSS�x���[a�ꕇ�0�;3nK=I�<�,�=��\�3b��E�F~_7���Ƚl�0E�.�3 ��@ �$�=�?� �Q���̗����4���g��=����*5��6�NNN�ςCJz���2@�O))���eY�L�F'&����	0������/Ʌϰ�¤BWr��'���xK��z#33�(�I��t��gar��J�3kqי&x����b��z<{���(�����s����\D����bcS��{K����S�&��]+ȟ�_ڎnE��k��P�,θ����;��њ�ݰ�i�J������W��bBFF@�FU2p۞�L�򺋌�>���-EEm�{���_^���/4����}tW-Ê;a3آ�39,Ǫܺ�$�Z����L��YpS��� �P�Q01[Ƀy��������ݼ	�*^�hZZM'̈<��`�>���i ��5�F
���R\�SanpK�A�@o���u66��f�����8��f���寮.�Q��0eeߠ �Q��ӳ2�Ī�0�B��Єf���o})�Г��[���OȒ���f�j��#4׈>���ɞd(c�@�iW|`.���?�����o��$S��I���!��]�kv�߷)�k��W��m{�85�pq�>ܬ�r�O�F������5Ë�`��5�����e�
�^���~C����tV/F��2���T,�)|�o1N��d�'�=���eb��T�}�xxb�v�v�u}y��a��CC���^Fﳌ��[���a����=���z P��{K��_gon5iC�o�������:i�*�Zr�'�RT Q|��������֋k���,���{(((~ ?�`uHR�).���B�]����9#���$R��#��`����\��|B||_Xゖ���_AC-�o[%������䖛/�V6PxQμ�)X ���&�E>.**j,�����|t�$���?ee�N�h��jf�B*K*�?δS%�(/�}Xk���e@�?���6Y���9cGgg�N�I�:`����T��;�@*�����O�Q�?�^vb]\^��+/W�wu�����n��?�m����W7
{�_�i�9_�+p�t�����7䔔H@��$kll|[�r'���J��,������geaE�íⱑ:ʧ����9�঍Jw$���+F E��03V��J����Ùbb� Hbz�&�220�L�O��1rp<��9(2gN��ǐ��405=8�1��|��)(D٧�a���3+���{����9>��(��:���:�7A�_��^d�G����};-�Ƞ�L[���Z��4�aȈ�~ E��b�e��X��iw~ #E�[1�y�T@"��\�4�;��|����Gy��)<cP,N�l���-$,�q{��K���p\.��3��=Y�W���� �a5��}���H�"��M1Of���`	�R���::3���L�l�g9,�)N_��
�?==ũ��9��"� �$�|�Z0�ِ�Tg���))�wx��P��`SJ��鏍�<K>���Q֎���������V���
��[��U�:�i�.��152�H������9�-mmwjj}cc�|���~yyٓ������� A���p�>>�򅨵%l�x�]�⽄t�)���4q0�������+�`<����ͦ�4+��{��,8f*M�x6�=��6��	[��,,8�����9��V33�5x��)k0�C#��M	��bRN��65g��NW��7��Q���MK;I &fº�W�>̐����.܁fϧ����DB������2yd1�]z�J�*j浸{K��Q�E�����x{�oޣ�y����uG�O>���Ϗ��xԀ�����}tw��xN����[%pt�Hdo*P�Ru:��?� F@�=TRR��R�G�-iB�>`��c�_�����ݟp�[��V39�$d?��j�Ǐo�OK�pR7��\@3�%ߚ0�8�i���Z@�΀I�?��j�e��KJ�:?��������������׍f}��ѮxN��la|o ��M&������y"��!�\FDd�{���Y6�C�nݺ���ްQ>��3n�B���`�E�:���s����QQx�M������]��_�G��H�'44�c6è�PQӖn���WK=��n��O�F������߳�p�T2�zW�G�Km���y�gF:B'd�N<��DGG707���Or�Lkp�+;���,�_m\pxDo��ͨSxt���V������w��3�յ�Y�?g1�	�${z��fO�3R���㟀faay��hy<�uM��.A����ߣ�_�$%q�O~x�Ⳍ��T�tt�620�E��7�O0ax>�ū���bt3����� '��W��Fh\'#��>q�u�kt���>���Pq7W����7W�C�ƙ�'������b����X���{w��?~\S["�p���Jv�h��P�22�أiS��;B�	��JV���۱�1���^G�������������y����|<^�i_��ߣ��f��3\��;9�(��R���q
K���w\k�Q �w����5@�5��O��G���@���Ǜ�@�}Ψgᭊ���epa�⻒��3g��>ž�0�_ҿ����u&��)b�����
��7�ô:����>������ʲ��w�7�s�ە+�NC7��g�� ,�Ӏw۳6$*�
gz~��F�9�4�ߵ�&F�O�XWCçצL����A�C �T9�.�u'>���K� �W�0z��i��N��Nܼy�OQ�==�x%�[���G�����vsfB�����*��KiO<�v[M-��P^�ŋմ���QP$Ŋ�ˀ[��/bb.��#�����m��F�Gɛ��Q�;��x�wr�x0�ș�����L��D f+�tz����[JՅ�*΃��n#mF��
���������x�@IɁ���'E��}��3'
h0@�"�����K9��5�y�?�e
�,�����2T�/M|c��_P�����:�[)/���$ޡ�?v��u`���^�8�Yi�"]�2����0+yec&���5��Uq�߭ZE�y���0 VVW�7S#��F	X���ba��C�Ǉذ

��_�Z0o~������J���e��=��7��oAף�]V�ஐ<�����Ks�htcڥy���%���4w�~�=���:ImP��	b��
��-�ʅ��D����i�E}N�U�;ser6x o�h�I�L�<%+�0�3*�����$�����>�{�e�%lI<���Yȥ?��@'�q����CEEE�QՉ�[�n���Y,�R,�N��xy-���`x�U<o����5$J�h:}�dEڃt���%)�������Aq�a��W���;��p�ѡ�.��o�̫���,��Ÿ���|��M@��r�Ν#GII_�9;� <8?==͟!���]�5WD�N�Qsbc�"</K$�*�*���p����쑗 צB�vt��y��:�<��A�s��Y$�W4`g��Vꡂ(U3M1�cU�Ց�_��::� ��i%�|Ͷ��@��A��^k@�p���Lǜ��;1To��g7 #r��8BN~3�{t�jy�#��F�lZ/N�I&�@��=\0hx�X)��T@�X�/#�7^�S�pummN�ӊ) L�/]�v�@0�f{���k�̸���s:"|��Y�W�G������\�R~B#��æ�䴅PT	�p��7�233�GlE����B"��wo'%%ŗ�S���oMQ��њ7fiiy��8q�<Kk�̌s�����ޅ���>��PQ��ZO�+��W�����[�Kvz��������8,�S�0����0�FFNN��\~�n5���]F�[�&$$�^|����
#�e�G�B���e�IIGlJ7�_����:�r�3f��&�xL�����r⁈!2O�[�Z��
�{jj,E�e��
��<i�wj��̇O$�~ ���\����=y���ӓ�����L�������jk߆���������W����" ��]/�7;P����-���$�����XiJ��!�k�LKG�lY�}>���yY�)��y�֝�G_��u��+��+kk'�U��;[�Ϭ"�tJ3���7��j̗����y4賢�?�����G&gf���5��������5�<Z���E�i/�-���x�(�9q��DHHH�u])`�S/�z�X![ۇ�c�g	e���y��χ��o��*+�;�TY)	�24OD��[x�0�Kb.�e�Qo�R�]���U���А!�/�/���䇳��U7^?�]60���KrzN��QX������{{��EE]4Դ�/��*q-�\|Y.�4ƻ׼ �q�23�?_y�,JE���l�����I�N��v����1*�3 ��c�q�Z��~�6������w�-�,����j5P�+Dv�8���$�U��˞C��\����;����
���
H	z�i����]}9��g�3�v�RlT��^$'T�׏O��>w���<, \��	�^щ`� ?��@popͧ��~?������J�~�WN���)����B?�������h7ңG������̲5���t <���쾅�+aH���L@J��ExE�]b��c�����9��	�4tx���׍�x7�B0Q���>�JS��U�����p�d�4s�������D�/k7�;8!�^MXw}��O����6=�u� �nS^���[Y�e]+�]I� �����>>g��&;s&���������p�D��`tIف��I��, �@c�s�Իk7�H���#l��c��X�N�ׯ�-�A@��[D��v .>a��?kzX����w��)��h�ÈD���U�g`��(���Ł��Q�E_�.���(�3�d7��@ò[7��@�1����>}z��x��ъO)5~�ZZօ�2^,��k9Tԁ^�� ULV����{38h 7��rsr��̏�sq��߶uɷ��R��1���b���xv���QŻ�#���W�q;����[����'��49��;�<{�{�����������:T
|] �5Cg`�RZZQ��e'Q'�n17~G�SU	q����[k������N��Wo<�s���_N��-��vvv�!��m%趽XC\
��P2(u���e��>V�$�x��ϯ��Sr ��$�ϒ���ů�ɘs����qל,Z�s�c�T��2�G$���bp�`�:0-ӱⴐ��i��A	}E@���a�Hw���}x��4���Ov/��ׯ�PN=�j�K.�������]J�5�U�s@ϟ��l^N����@b��p�X�3�4�G N\��?"##�}i۰��Ύ7�q/'�� c�ǯ� ^+O�@�86]=ѕm�wcs=������*�~�vu��Š����U����.��*�A��>����b�)���u��S]-ϐ��=� !�`<�g<z}~k�`^�׭�6�mڨ*��3�J._�7�U�9�~����胧[��k��~�赓&��?�|g��ן�E���a�'4��wl�ə?>Z3��$0��s;N�Ol�}�.��qh��9q��Y�	�8�;�?C���(��+Y��L=1�T�\<�_��s�f&���-����[l=��#�;%e�������2�#����ܤ�K9��A�Trn{�T������0a���&3�6�g7R݂��\�l�����P�sss	s\�Q��b���F��|�	�N~��ܖ��g�";5�r!�=�HEs4Z5��<�(����4��6J)ݚ�ߎx!a�G���wN�[O�b8��g8�0�,&�J!���"䬟����#�q�7�V�jKO�$���
K ��換5I5���&�=�a���
��
b.TP���(��0)A�t�ۧ��N&�JT�9 ^/Hɢ0'o�M��0�h������G�[����%B�V]g-;2�FY.%zś��0�zW��'T4�]
B}�{�5��p��R�Q�l�w!�t�3Clp×&���{����-�]ى_r՟롨����W�Cf�]s<|6:W�pq[El��8)�D��@�2O%L}�I7�T����J�x�9�ð�Aq>�PՐ�z��h��φ���N����R���+�!�>z����5�dU�R���<z��r���Ũ$�r%����s���k0�|kz}�U�����Us8���?���n��5h=3e�������	�E}�koG%�\18���v�N]G]�"�v7|g[��Z>����ZPXX(��0F���b�09�b��Ѐ_��WF�
��~|b�>(�&]˳줲'���:���imtV�o4x�j�b�'b_�<Hvy@������M����C���ש��o�K��q�sa�0����l���῍qb�0A��bz��y���Kn�)_��;94}�O^=ejfv�-]�{�Q�>�/[�<=���������u���ى2^L~`�Վ�׆O}��.�J�Bu[Uǉ�ʊ�&E��rғ����]C��'�/!��r�PꠝIIN���q�,s����İ�_V�_IMM�(qYmj�!%!��0�3�8R4�c�ͫC
�dW��-Q.���&��	����Q�>�*��(���o�wHuuu�J:���J0�[U�O=�����Gp�g�s��H�:��a~�g|�GEp�|��l{�T� Xqjݖ��ۍ,,�X�i�+)��'ZP�:�����K���c��2;�<m
z��yx��$�=o�۔�v�R�JR���V��V�z���y���X*�c�g�u�o/�T��r����x�ncy6^�����*膭���||�_v ��&�Q5:�0 0P7n![J��7�t�@�'E}�:��SO�x�lo�qrr�sE�Q0��e�)=~z�a`�pL�]��ė#�P~N���� ���ts��uN �M����d�t���Yv�Z�~a5[mS���'U&�����w��"~kd�צ���-¢u@���S�\*���#�)��v�����k��Ӟ��Q�\6�ҋ�ذ0�,�`M9�q?P�B�夠��^O�|Y7	��?�-���6�o5e���W��o�Y�ڡQ�I�}���9�"'�z�'�����OA����*P!Zp,����T�l�H�=|��X�Jje8�����fGN� �X�
L�N�ȅֿH/9�L"�z�F|SZׅp(�3S��yx7��7.�L����疔$[л�2�;��V`���qP�lt� ?l���Mb�*�>�����,��_~n���\�na�\����D�U�q�F�9,K�t^��]5���Qg��|�N���/�	ص�f��?�<0��L¾�IZ�/J݃��+A���0w�mW�����J��J�b��	�2��wK���d��4K;(�8���X1N����3�CY�EHM%[�C��h���%���<�ȡ��}9�>a�Ϧ��*��KL���cϊ���b�dA�&����o���bu�� ƛ��tt�V�C����;�Ď.ᕈ��[i#�GƲ#K�f�|7�"�LIѻ\��Jr"�"B���u;�s')��|��m������k��-��a:�tU۔��
zB'wӠ��9>w���V.�(v�|24!�>�"�cg�r��"�8�I߱�-���a�z*����'�w��(izgf0x�=qnK�:,�s��� ��� ڿ~�{��k���9�h���J��^x{�/�г;]��c��"
)��C����ߡ�÷ 97Wa��#f����|q.ө�4�©�)z��&{����K�
�U�J|�9A_\ �@�����jy�aG4����S�a&�ƻi֎J��_��Ѷ)��������8�6�_����ɳ��bތj�P5d|xt7��\p�X�U�T�iS�΃�Q�tH�@��<��")F,9ӥ\' �Y��8�m�!Z�(y���8֏�E��9'�BCC#;\m^�(�G�`\��互�E}ܳ3�+�I���g*f���ޤ[`ݗ�B�~%첂kS��l�棹V%�J�D���xc'�,׬���s��{d!0YC��.@��h!�7�u�q�h��x�0kS��O�}��5Rh��?�asqǋ��3�� �#rmsO�$Œ?�vd��pi7�P0��z�\|ra�2�p���݅f��@���/���-��q���|�u��/k�،�z��y�B�a��V���o�_ YD	���	a^>�@�1tbG��߶�ڐ�k6j�R����Z����~cbx�6��c-������l��p���|?��״0S��qK*���%�����o���ڙ�β���mߒKd'|k:)H��j��WI^����ڀ��#�_�;Z����s/�m�e+I<w�{�K�W��0����T3nMVP�َ�v���y���eS�����+Sr�_�'P�[�̍f	�(��z녝Eə�E�ℍ&���t�RL��T���_w{a�]uI^5Q��/qy
�IO0��#Rv�h�Z���=�{u�On>rr�G1Eu�n�>����b�jޚ���6>�0H�m�JX�Є�Rh| b=���^#A��ps����*\&��@i�˞vY�`ѥ���g�s�7�Q���Ű�q�N�������޿�{� ʝ�6��ٟ�|&�>��1� �b��j����0��\���f��'�C*՞���,���'��#�H���/Z[s�v�=� ?dw�:���6�S	�nd��5%>,ՁΆ�J����G�����YO���8�ZbB��d��.]��QN'{gD�m���	�2�r@�D�+c;�J����x,��2���|rJ@�� `YOT� �o�2�&cR�w��BT�[�βz-����Z��`f�ĉ�8%�1c�;3��z���%�g�k6��F�~|�h�Ҕ&�4ǞN���|�7�s��-����?���w����Y���Й�I��,g���桲@c�:88 ��X�Я���?��c �qܗ�d���޵�W�̄W@ L5$�~�2'Ǧ��f2+�
����]*Ы�<��$Y�;Ѕ��,�*�**��� ``�A���������~�wha���{/���~�mݓ0O���b����T��,8�Z�y����M��F�J��6��8��Y�| ��'W�.p#�P���� ��8�W���c��
���%6�l�N�����z?7_S���HlJؠ�8-���3li�+D0�'5��3K_@�V�*���z��gӶ<�C�/�pjJ�ʛ�D�U�*�OJ� ������>M;�:�.z[��֦��v���b�= 8����w0���FF�~	���:�o�"�{S�^��Xezݙo��$�)0����܈�h��W���>���f�x�T��
ֵ$�&��ѓ'OB������Y��5���n:��y[6H� LD�b����_eA�j�zw�N��&����TTT�S)�A��_���<` ��y���0�rz�7O��4�,֧�8���f��{��J�-�?�2��:R�7�̫��u�����~f!�3.z�E�v��20�i"*}������ Zi'i=^Ì`��ۡ�*�y. f'<��B������>k@����J�.Jd�(����lÊ�ߛ�������>@<��g]0s�����[]]`�];.����Tc����y��*��B���]�(�U�D6�qI��j�%��B��w{���л�@h�t'~l����+:)�8ۓGLF��wx�H�`t��%�ĤC��Bo���g���ѻ�d��vI���<��B�de[��32�����Z]Z{�z�!��ov��/L�X�s-��{�'E��������fyӎ[}���������2Ӎ+ێx'"(H���T���^�u��.�IzW���1jkM%R�Cw��X�oi}0wV��Ӳ�;���eid||Sq��	Oqo~9���k��ޖ��?߲��%�|Nlz��:���&mb@r�tp�%�����]t�̜&��!;=LrZ�e564�0C�x��t�C���w�`�K=��W9�_�&��i�1�;W��N>���*��#���86,���@4�2���|;&��4-�**��T��g�k�HN�H%���Ͱ#���C�|�'Kh FOenqV72�!���cr�����y7Y����,�ł�%N�)��s�*��]���U��s�i��7/��h=��U�$��+ը�$v �I�d�um�ީ�ק�0�~�3���S^Ϯ�l�eZbG+��˵L��Z�wU�!�[P���	�;�C4g����|CF���44�w��A�o=/ۏ޽t��'�wB�@�����Z���R�E"���buWН��%��=w��GReYǳ���&ZO��U�Ӱ/���R�G�� (�M����,�h����e��Id�KI���ϟ�2�D;��������8&�n�%�U�~m�;�i��e�箻��IHԛ��Î��0�=�ĕK���f⫀�u+o��Qٟ?�C�}:\�+l;x��3����O�����t��$vRn�*�N��贒��u�諠:����땩��9�y�%�w"��|�✓ghV4Bf�Om�-��+��m%6%�<y�w���B�zgaB���&�l��ڬ�4�3�(��m�0˜a����� ZvR�����h���Ԍ����`D�LH^2w���Wv	�N�z���s"������maI�j�~p��K*��y�R���K�x��=����k�i{,{�y�t�Qז7�Ӳ*�۔�������Մ>e��S̭к>.T�:z��cr7Ȯ�8v�A�0S+������z���}ZЌ�d�&������)�z���K,h���V����=�ǯ0RF��@E�v9�S� '���#cc�N���?�@�jU&�ge$����XM��B;1�x
����F�` S
�d�������У<2!�x�6�ٲ�jހ�0���uAo��?��d��p��a�?�hHUM1"�wLj/��������<���n\ȓ(3�ԓ*w��⬮��m�ȳ�=T!Ǳō��j^l�뙟��Epx��Ę�D���`n�:&�
�g�S��ZxJٚq����`�r�GM�VCB�f8d7�0���+�P��ۣ2�l����L��d:��QU�a0�N��Ī`�;�T��<�kW�0�l�3�7��{'|٪�����)��<�o6P���s�v`W_�	��1)���X�Ģ��7������J\�}�F��er���r1�-�G����8�<vQ���V�5@'���2z�RO�L\�s��@O��Er&u�2�ޣ����RO4�r ���ׅ��ݼ׀D�-���פ�M��8��ʙTگ2�-"q4U�؉��->?�HC	��]���;F4v��럍�Ր�
�3� �yx��h܈�&s�X$��+��?�����Up.s� -� �C7�50?�[��M��� #H�o��s�,gd�2� H�BV3M7����b'F��Z7П"��F���E�<?_S#��M��Ĭ��L�D&@d�+c ���tͰ�/��*� ��͋��)5Jݷ�����ˉs�/�rfh8�s�ıQG�Jjev��iZ.���\\���=��<:����$C�_om1(<vkԵ�nzX�tb���2!��٘`Z�ߤ�&��"��	�{*W>�C���"/[8Yv�΄W�u�q�קUT9eBt�N表a>[��j���&$�ͯ��L�z�/¬Y,�R-�p)�ۂ�mʽ0�]�)R�"�����w�Jm����vy�������M��u�j�F���L���0�\�62bdae5vsMNNfd4�!��P�Uo>W�f;J
h=D]�>����+|���0��;:���:>����af��}��ݲadK�
Z	4u����:W?�أZ���%�&J������Sh�RQ��J��V��1b M$��o}(�O���D�?�Td����"1����f)�^1�B�*���x ��̵w�l��zL�/%<�B�\J��I"��io%�/̙�l�	�";��^M�	?�ۆ,ŷ�|C
�dXNl"ͦ�!�_�编s��/�ښMlFcr�m�L-�~I�r#߲s#�~����V&1���0G����IҼt�qR�
(�{�_,3$�?���J���!��sJCN.���8�ķ����1r�u^��m�*J?�WQ��ϟϚG��prr>�*MdAW���U?�V��tU�_kq�ˍlܫ����'uA�����0���M���?�
����P�^�]�n<���K�eέ����Ji~�PK�	q=#CB���a���s���'k��*t���=�zcc��T�[��|UUU�˚1������S@D�*V�e��&���E��u�k_K�J����414���4��t��ݡ� ������ӌ'���^uRi�uy���/����"�L5��Y�2Z7���bB8GG��>#��t~T)UӬ��xx��c��.�'1ܠ�	'�4�dhw�Ǐ�����<�i�UX%��?>1F�/�у�Q:�j��<w��SR�.
�����FƫW�&WW:�X-�������ǩFa�lm�/��$`�9��J�c�6����j'/Ͻ<����ʦW]����gs�,535��k�&{��l���̀��xM��5pĹv�!s��6�ȥ���=π�  @AA��i��5x�3��
�0��J}q���u���L=�g�
	�o�X:����㧄���|��H��>�@��3�o7:�����/�]���#:<�lO\�_S��,K	49L�|'$"(>X�q���@{̈́0��S�w��^^u[��0����O����h��~D
#&��j�W)�	�I̸�`��Rb��-222�EG�(ˏ�ٺC�A�e*�n���m�q�V��:�Ϲ?c_���2��*G<�s��Z���u��~a9�n��`�'?� �~&����s-�%���cgJX .��ci���U�O�ǀ�]�2�<�������_-�z��q������=#�LS7��΢���k�L��Z�w7�^�4L �wEF�u�j�����ELz��L�_-c���g �فzGLP�$�XH�-�	�R0�|�[.g�~�!�pa��ؚ8M��s����Ǣ��d����!���B��[���P
�+�}o�w�Z��QQQ]��]��cG��넳��񰳝l(��n�T���^�m�����*�9���p_�^�˚�b\�s�M�5�/X{:���퓹`4���>2�C��F��OT�bn�a���lԳ���)�а�俱��Γ'OF���
k�p����FD��e���8fMq�@E��aZ���5/�;��,cZ���֭, >3Z=S�OI]��( +
h�(f�(��/�8Tl 3�G��^);p�����ͳܞo8䄈{I �.�@:Cy��-�6�c���q_i���M�{J�����
��'�<[��@<f.��8���6�φVE��l9Eqzn��qs~1�������Vj9Į(n�%��4���r4@F��ss��"�ēkz.�:̾���_GD����v�(̩~C~��n^�f`��W��L��+1R�kߪ:�M��
�p��_��W�d���/��F� �nA�ToѢ�>����l��[//����\9�Ǵ�C�� ��.%z�K�Sӝ�p�?�J��9��N�6�6��F��Lh9Wp�y�e
O�����f�>���l�����$%o��r�UHڰ��߿�X��P�m�^"Ƙ�m5������p����&��+!NSy�+r6����{�սc�a�����"�����t�N����1%�̱c<����W�_� J	u�h.q�	�lS���o�����Jn~�/ej�7���&�eN�F���, ��m.f�p��ۗ3�8���nC'h Zfj��G��v�Y�����'����=���a��pW�׽���K"�`r��'My[Rne0��,�����X���B��qZ�M��ڔDv��=��	�H�Z��p7g'nP\D$�9X�9��!�C9�����E]�Ѽ���n���j�N����AP���l��H0��Zt�(��M?���[b�s�[�8�Z�z�\�3�WƵ��O1v�O2��[C����R��z,�Dq�W�^//QK{��skCj�Xw;[n��?��*��ɶ�|��vG�prd�_�uSu�$䭽A�g�9�g-�͓�t�=��;~k�,N@;��8n�8��N�M�Ra2������IJ<��ȾbA�����  8�N���b�E��~�F��v�0��Q"��Bk=T("	��_�>H� }��݁B������@�g2��0��(a��c���|���+��ߘ�v��tuT������ּt�E;�.� ��w0
��z�4�Du۽��e��\��� �"���,YVY��^+��$&to�ILꯗ�%�t����vG@S�\��_�}�.wwq��ͬ.�ż�9�3�9"�s�e�L(3��֛=�N������q1J��0@;?��+���-\�C�DQ�ݥ��:�xh� ��h�E��
�+�����ʉ�>�2�f��"��P@�酲��7��-��c���?����ܻ��?�y�ϼ���Î4g���KD1���]��o��uw��� n�OC@���9�rjr=:���3v�)jP/S�N1=��DO�#��W!N���kV����+a��b���w�Eo)�j�����#��B�3������{��,�����l��#�$4�A�
|)zr 7a#L.�U��W'~�bS��y���S6�gS��0ܹ��hl[���W�bZ�������Dsg������Ho���:�`o@��z�%yYW�Pl��ֻ��D699Q����.�WA`�sj�<d�} ����B+)*�j�3� ��i�� X�ej������ϟ�8{P�h2��ӧ�D�UUG
��k�V�q%��t��d�����@��Ϸ�i��H�{@���u�)~���׀>�Ud%.iCf/�D�_���� ʢE���3�y�7��!ڤp��y0�~ �ͯ�$����{�:��J��-�'��7�q�A	���v�^�������]:v�I�<�徫:��:>d�;�4�h�� ���;2'ɴ�O�~ �e8��?:�Sy|�����	�_&��VV�LШp)b�,�ߏ���i��@`o���qz��4� ] ?#�,��l��
6�X���G�D��R|{w�R�C:��׮����w\ ܁����ֳ+T��;�� L2s� X�f^I��0)04�8�?]�/^
�6	��~{�
�q�������&�>���$�O5�E]��!\��8ا�=z����<_Z�ey[%�Xq�}YW'��8̠J�z�J�*�/�z�2{�y�cW�����c�m���=���x�U<�"��3ʄȻ������_[�2��X���2JN��/ԋ`������R�`�W��b��X��U*\W���)�s{%�%���O޵D��K	p�Gā��h�wj��������h�̐����7-�Sv �ݓ�fP�lj2ӊ7�1�Dk *ꃉ�o��fy.*��)3 ����𖁆Îl�h�yY[Qq�g�˛Q�⼼o��ӟ�1/聚�95+�����M˜��T�{�>���/�Ҿ����� 	� S)/�.Ɵ5,Cߗֿ�����oa(#	T.�4��ud�����O����pо~�����O�<S�<�~�u��!���47R��eؓ��z�������$��%������E���d�2�:��ս�o��SRR�x�lD���~��unJ?�j�;V�&�g[d`��Roh�!��f#��j�? F���E�>��g��N˻~���)b�Ɔ�;[��Ӄ��_�%u��n"��'6��H_Pb.3��hY�m���6Ϛ�DKI�2= �e����c���_N����S�D릜�mQ���A�i����K���M�>h�<���S�3oW'$�-�}�9�ϱ�	w�{a�R�e�|�] ���H�}=W$_�~��2��'�U?b;�L�4�ID&�E2�9���⭛E��קi�%��Ǔ0q<*y1�����|V�y��~ˮ�ﴥ�Fv���x!�
V�X
�쀇o��tL�yl��;�؈9/��X����HԢ+�:Q
 ���!���Ͷ���|��#��\, ��h����Sn������&Os*Q�:��i�]�o��5A��yÕ��o2��/�R��Vi�s�q=��	�7���[��D�y�i<�@\F�����=8��\& ą`�hF�8�1E�R�2u<C+/m�X��K�����	�nY��l�5[`v�8��Z�G��0V���t��MԜ��_d�N(�:�Kh�?��'~�0^{;��������s����mÜ <�
��̰�'|��iU[4�oI�}����M�-�YK}�@Z!=�Sx4�m�v���ٸr��r05�>ѭg�
�O������E0ЊZ�}�B���U�k�8�㹑F#l����π^�"�egr�"�l�	hY��6�!�wn��yc!ŏʩ�^�����@$p#n��0���O��[��=X�([� ���ǕR�m!���J�6<D��Y�Z���`f�R��td�9�p��	r�>dl�q�8��������n�V����}Q�AKK���!j��kj���٥mx�޾kQ�+�_}�I���XI]��N�#�gNsU*eF����FiC��u��£��jr�Q�+lǈ���E��h�"�WMAp���@�amb�z,�.�O?<KCgh����	�d�1g]�vm<Pb���Ṋ<���(Nη�^*CM���X$������޷��###�a>G�\z?O�)3�AgUx������- �N�#y4���3��8����p[�52���/ý���H�j�nɢ�\b�<�G"�\�9WF�*c��Y�ѩ��ʃ��b�zڦ���������jÉ��w������/�ȫб���Z�I�up#��_C<�u�����Ҵ�z��6k�低Ӭ!U���廱�~q�����z�Oc�ŗ�m���(���0�N�� 3񀁧���}�ŵ�R�)V�y�&-L�m8�i������$*&& ;;�ŰO����R@}�]w��İ�N
�n��]�cw�d,Wl��5�v��s�+�?N��������)�Ua^���{�� %��ςx`�W�ZM��}HTԏ��\3Pr[O���S���U11�0Y�nl+?�/�@x,y���-� ߨ��鰩jN���'������eǭ�g+KO�
7PR���n�����J�g-���Q�45��6˱��t��Wa���RϞ#ܟ��������>UX�gEv�W� X�:aH��a���`	~c">x`=p�g�&�ڞ> �	�:�-��A�\��Na����S՟=vsF�<[�-,:=��6A%�az���Gc2����&<'<�ޮ��_{߲W,�&���շ����|4���*�cy���t#�f�g��/�x�8�z���_���� �'�###?�-��Y���l�jP;=�*�v<�̓}oA'�
���@ᕣ��$,�VGR%� ���s�����a��5��0��>�q��5�7�M@p�D�~Q_�cTXZ�l5<`X�Z]Q����Qv�a�wx^g�?�qg��b�+s�A-`hE�z����j@d�����j@񫘣���]E�wov��Y3�Ȏ����XJ3�U�>O��;W����f{��uZ-��x�bn��s�z(u[�n���^hom��̶HBMd����J�ho/�m%�}vp*N+�*44�p��>����\���F�egV �5���c �v��U����앬yQ�{܄�-����M���9d������P�òFgi>4�\���������B�a浄�[SG��jH��k�\�3�=����>:~�ؿ�g_x��ׇt\M�{ژ�I��7(�IQ܉S�X�m��p�.���ھBEM=�I?3��m���;F�)���q="�~�ds~(OB7��~O����@�Lu�����XZ���w����*�T���`[x������g��n���:9 d�6�3Pj�'}��R;<g�KXhH�_�pE>�HT��/��Y�1
�����Ij�؋��5A,VP��Àv"�g��Z��B�7����>��tv����I��5)]����hZD��	�^����[�j��%o0u0�䩿���v�N�+�?.��?�xý7P�\�%�ݳ�)W]�D��>��I�*�miQyg"�˕�J�B���N�t��UfN�gI�$�5 D��p�K0����ik��f��l����nG�eq�1�-��)-3�i�q%�..ش��׽*�fS��k*+%j۞�NO[d�Pd��$�
���.�MU��)�5]A�j����9���}��h�1�=�k�}˘Bm$�W&��Y��4�%n������Ş��v	���{��m����}=�}��b`��g<H�e@�[�JU�M\)q�Tv�s�N;�k"{J��>d��v��vw�qY���*a��v�;Vwm������Hk�1�5����z��&������Sy�;%zK�(�f�~�遣w��y,6�����وT�줹g;J��R����'6?x�^1%w,%�쑡῵�����>�.K��K�Y��`�g��[��:�#V�Iɕ��'�\�8����466���-�����ǖ5r^,�,�����b���K=t5g�j���E��`~c�	��}\\��O�� ��>����1����m�.�ˉ�����6�1V�%�����PP�V&,Y�()	� ���@r�Ֆ55�=p}����$ҥ��>ǧQ=rZh.�����	�lѾ�	8�d�+g�����O^^������!9ᐨ�ҥ�똂�����:���������[����WR�dk���tt�)�-���g��T��[�e����c����$~I)^OAl$D!P`$�ұ�Oh��r�%Ay9sO/_��(���ﺪYrr ݛg��M$]��t�:?f�oĻ1�	����+��K�z.x·��t��J�Q9��=�ug��;�H�`��W]�ex,������U@�*ym��x�?qu�Ǖ�m��rk�ߙ���i�Ef<~2�꿸R�`gjε}�fo6� �J���pWl"��ʪ���[`.�����������c]��[��	_�@:�b�8���)�2������}��7���^��(��_�ԉUN?��ݍ].���o9�����,u+��5��8���ֳ�6�͎O�y%Z}���]S���H�^�����n�ߛ#��ʔ���p?�8�_�X����]��8w��JJ'�H<���bѼ������\�%N�X��. �>>9�E�T'���\���ԍ������U��lZ^����Pq��$�/�_�F������͟��ܹ<pb5Fi�.�7jV�j0��\$/bRp��ĝ)\M����Ϋ&K����@� ku���>jqā���.�NCj�:����f�ڣ��wK	�����+)���w�b�4t=�|�|	C�z�#�m���w���=� ������T1\��B�{��T"��	/0���Jb$z��������]D=�����ew�0�O��!�p���/<W�=L������0�+�,���/���=j?;�ů�NcCÛ�3���NN � ů���4}�ۏ�����<'7wr��{"_׵LK�M���Kx����}:���R"l7,�����'�m�*�.ۚ���7wM��N�}�����Y��`Gg��ҁO����|��m���9�_=r����o7\�;�,JM!��-��� �b��=b�(vd�c�]8��и+vĀ����E��m�� a�4��K�i����W��k��� ݾ=ؘ/��s;IzDb�OM�R���>#'W7�q`�o	 n�z�������f����e|{<��N���{������;������8E=|�U߃�\�m�6N�$��TU�}�h,��n�-^��9����c��}}�����v��Ս��ȑ�!�& ��^_��Ғ#5�lW!�5n�T㹘=Ak����m!ͱ��������
�~��= ��[����y�`��|7�zc]I��3?���������k�ց���u�,�O�����B�b��J�+k��W�����}u{_Չ`�ǹ��9��s=C0�r2�.8*�P����O�w��O����z���*s� 50����H]�<�Y/�o����_|k�ؚVŃ)��J�.�M�瑉i��`0����`��x3TC�.8ܪ�c趙.�b9t�м?��l��jC[��}�CQsppLH�t�y�����Ħ_�x
υr�	֑�D��vR��_:�9����~*x��W��*+˯����g��f��>פּ��'���͆'�k��:�{Q�*%���U==ZYY՛� ��lS>C�櫷\����i��o���ڵ
�����
�K�w�����k��K����!;?�
��T���'+��V�[
�xܷ���-���HƵ��|ll�@��H`�H�O*��z���}�ug��V��D���uuu	���*M�O��r����M����ƪ�����ش35��1VG����d�f�B8�[}�~�F-Q�%��FwNCG3�*l��o�f��T����������*2ɍ;���<	��6��=Pҹ�s���Ͽ�/�xɞ�k����}{���Tz��U��*����62���eQ@+��Tھ�W����i�	B)��Fϣ�yt�bLɍ��eɸ	e�;ӿw޴m?dZk�̄ĀVC+�R��둂�0��PY�p�Nccc&AAA��4'@iR�|�aW�㱐%�n�9�ԅ�?��jFB�9��jd�̤ȝU��]lKMr��pX\�uX��53*��:z�<�1�k�I��"T���/�5��+�����#��Qe\j��G�u�S����RJE��(��M%3��)$[��TB6Gvv��8V�N'��8��>2Y�������;��^�^�����w~>����Ox#�����st|��ق�"9n;w�g����{s�=�q$gW:�N.o �q�GJ�_��Rg��<��t��S�x���*B��׾���M-J�K6�o���=����u����q��U�Z���h��u�M���h���2�j���J�vފ$�R���Pq���  �66�#˕�#lD��=��m�%��"�frQJ��x{�l�eE��c����;/�t)���4��r\�{�"n��D��`5�(��wWfo^(%���ѕN�MQ��+�g���YYY���e��a��OMC�������[����&�������K�h����^I�+����OVS=ބ�_Fߤh�	A���ܠ������+C���I�t	��#�0v����M�=���bEA^�^��?>�M��O��q��f@�L�&p�.<�x�M���gV9�j���Z�_�	L	��uH�.v�����^���~����Ǽݺ�J��Ȟ���8��~k�-�Uq`z���˅Zy-KK6��G�\����XM2�<�Zyc��K���n�ߩ�;99����%��ݪUSwp�C��}(D`FQMt��؃�&'���Ϸ q�W�V#��jܻlwoOj�6�	�"0�VǑ"Vp�s�Ǿ��F!�Q���;Q�� �����E�6T���E?Ju�(U�fXŷy������l���}�S�8�ھ��+�ۛ^�!�H5$�lR�/�"��<�/^�p��s#��(�<^p����77��m�۴�]��y����e�Sn��{�a-t� �3�{�����#�}i�.�xЃX7���[�Y	��:xe\Dcs��(Ɯg���&l�Y���{�{}U-��&�������T̹=O��P�^�5h#��}?`�������#��n���nC�������c�����K?wZ���\w�m�:��<��
��p+\9�~�ɀ��ɾ>s����g�{*���o�á��C.�/��&��_PF�D^
e����UI*{鮛��uW��~Xhl�wj����u�Z�B��Ab��aW����R�*$��.\]}�t��;�q>>r���֎Z��s�f�?y��2뾽����זֵ�!IJLE�yP�:�ء�\{��R�*�7 �����MHP�0տ�������x�'�1ٗg�<�3uԖ���6�Y�?ˠ���ɻ��'�Bw/��6���v_��Ʉh�;T���W ���)$D	�ܓ����@��cd/��)�з�`�������Ej��SN:�W�l�ΐm6`�p����q_�MZ�����.OwY���Ð"ᕮ���'.4p�K6�-L�e,�~�5]����9"$ ��C�5��b{p�,0tL�E�[.B���oH�С,���VV׏�Ԅ�cM�?�U�������=?�w0K�ų�m?��p��6�� �$�CӬ���4���\�#�z���ԺI�?�}ܪ�ېF��}���<&��C1y�ϽA��V��T���O^��@�)75�*���+�"%p��	��/���虼0�+�'�k�(
�*�~�%(�o��ж�Ѻ��h�'�Ȳ��hr?�+Y�y��ၰ�\��1��0��������`K}�҂	d�|��!�)C7C��6J���g�C�ʙ�����˵ �����x/�ؿs,M�X6<�.R�O���$/a��Q]��<��}�as��µ&�HHZe��EM���2;�.��U:�zFֲ�߬�Q{Dz~����݋k��p�Zԉj���Qu�А �|��7�Q�n->�%�j�ͯ������Z��S��������!�����������Hf�ɡ��
��rB���QH	�TF٬��K�6��D{M�_�'a�9�y���e��9X�̎��
�^�+��X���:= $��$'��vo�^�z3���\���ׯAjI=�BcD4����?�X[7�g��:�M�y,޵n�E;'�X���f�pOY��z1���lF��q�Ĥ��G��KJ�z��]��y>�z*���7u A��FQzq�s� �Ǔ&�i*$�)ڌHC�]\�sc�'Ap������D�Λڐ̒lH���͛�%&�����V0����j�ޅ��>��'�Uҹ�
���$��J����A�R�.��5 ����O����^m����??��6X�~1�+�0ul�ʢ���`bZ.���^`�L��]�RN�cy0�q��2	��R��Mi)��� ���U���Ь����>��-4N�5��F���8y������D�L�$i����e�d���5�ى����7���Ŀ�=!�I���=E����W4��ʨ��H�����⍯���Y*#�z.+I�>�߁K����N|���Y��X܄�\��#������n���i.S�|%֥���7d�f3���ms7�K�~�c�����osA%��ٰ%E�P& 7h7X��+#Z^a����e�<�����~dM?����5��r=����BV�D�߁M,�+Xӟ��!/+
-%iIl�ȳ�S���29�O�W������˚x�>�L "" ��a���D`��q�x��l0'�r����:IL�rS�2���>W�� 
��3ȶV�S=���C���P�l�ϻ)c:�R��P���������b<�S<o� �
�� �'������2�Yvߥ���2Jm>x�����$��)�3N��T�;`�˦�	 ���.�;�OBsR�Y�/\��.��UGu�s�`S�vE���,2�?b(۟ˈ��ʢ=?����K9��:P���)&7�$�oJ�T��[� �yzz��ᘹ ;��C���d��R*FF.����p+���Կ�tz�x�`��|�� �o�Ѕfs�p�T�޺ ���i�����\bp�V����K��ڎ�o�y��ҳ#��������0.R�?~�a�����ɤ���>��O�dR�[����Ʈ!��.5+�_�|�	�*q��]����?^;~�.jL�6/������U��Ⴂ�囷���1�P:�57
�ef��Z�Lp�����N�o��1-�Dq%��ln���Pd�S��ı~���7y`�,T�_��n�,�*מ��-:n��%iS����z|+ 	��1��_���gil(6���7�.�k� ��T���o\��Y���q�l�rp�*Ɇ
S�H�JuF[�ϼdl��*�n�] ��a�.B�8�[=
I��V��*�Ĕ�e�}}���@���,
�!�W�@ZF&f�+u��BɃӣ�>��U^8���ZN��̆���
�����k#��ɕ8]�����6:�˨�N�о^,j�$��쵵�>�LLP�2%�-՛::�}:Rn��-�^ݟ0c�X�L� �]7󳃰�'�X�����$��#� �kTa���@��掱��g�գ3\���0)�����j��TU
.y�K��Mz�h8�����tX8gW�5ԣ�V�h��V��e�{�~(��lt�e���y>kzGl�L���������,U �tf�f�����&�� Uo&8.83r<M��`6^.��n{,�iO��a_C#�B���U��ك���߮߭�>��(����5~P�������\����_�Y�
`�3H�ٸ=��"ָ.�:X��2�;�L��/�!�����|�ϼ\\m���lU�N�oũ��{h|�i<^�u|a�7ċ�zmkۏd&�{����ڏ��7����6�bc�a ޯ���p�W�ߪ�$]s�ĥ�A���C���nt�2O-n�kj�kE�8��L;�Ⱦ�|]c�1�c�]{��۪t_OO�l����q}|�M���G	���*º�5cIFI�D/6nY7�=[U�;<��"��}�!�8��^2�g� /ǞM�~�=A��Zo�׈�J�9\��TV:�<��j�+��i:4�4�>�r��8�.�*�0�d��u7e?}.��B����qG���l����ɖ��;ގZN����2Ӎǃ'�	��5�b�ԑ���s_�O��m��[X$
��I݉n|�NY�D"�h�~�����Ǎ�@��O~��7��]�����2z}�>S���Zك����]���[�(�������A��
��Ƙzz�bkfS�Gg%�����-?�F����	�@�:�=��*�������<Xo����\D����4J�5�o)� �6X��t���\���-$}�סNZ��Ĵ�ѣG�+�1�T�srS�?���/\��6?XS����3��uUA4E���ۆ0��澖ϼt���h�.�\Sk�
�=:��)z��6�ֻCm�P��LJ�f8Vp������:ɡ�M��M]����c<�Ht�|��P)�3Î���>�q7��c�\��y`Ԛ�T�.�t��=���ω��V��x|q~R��c,R��,?I��vee��Azl<ӎu�J�Q�_�(DX~�y,�h�>EG-f��C]�cЙiЧ~պ=�L�Pxl�����@N"�ߴ��{���TY���%�"ή�/�}�}!����"���\�>xn�B�SRP@g�7L��A�:�r�|[i<^�����Y�<��ή�hVj��Ɇ����s����s����6X��"��˂���Z G1FA���A_�m,�={�U�j�}v��r7�qo{��m�+T%��W��ؙ_�߆���e�=�*><;�g�u��b������,2�˺ꆻ=�q:�����8J��xe�x��D#�W,LF"0�K`�]�+tR����������?�L�b�g̳�]��_�F���
Y9��9z�в��.Þ힄���6����Y��.)O�xg��;`>d��&..+���ee��8\\��ν+�ԟ����27�Z�<���ZZ��]�3�w3q"�)���	$���3x{��Dئ��m�T�v�����KLBL�]n:o݀���o�h��ң���ߖ]M}|ꋎ&�wl*�.���,���}��:������h�S�ǥ4����R{�!]Z�&�ΐ._E���&�!�y"��	[\�q�)�pCx�����A��Q6�Q,�`�.W�����B����J>��^�{}*�|������
l�ΓC]���T]�;L-�Cd�D��B��\
Ŭ��cR�e�;m��]�S%\O��8���N��+��oۀ���=�S����YiI�Eǖ]��D��/���QV6�Q2���Q{S��^FF)���{oJ��E8t��C�2��Rgq�w��OZ�7��i�� 0/0�����הL����6�j�U{��'��w������(^D7�{���%��1��'��m=�ZMPL��C뜫F`���V��ޯ-�v�`��8:m����J{,d3��P����c�J�p��.����k6�U�_���ݗT9���y~�B ^�C�+��zx��2���t��2N�4I��r�6�|��ڹ�������V�<Pι�QNy�N�e��@Z�yF��,����mt�)0	6���f8��	���p}��v�#��d7��J��+����#]�(���{����˭�$!4'F��wm�"_~tSi�'$_���}���C'w�ax���ϥ�C�����y�~��!��������~]�H^�6�����`[W��O�ݫж�l�����`\*Z�+�DÙ��M~i��2Sv��)3�����<�g�?w:�s��ﷰ�� 'K�)$��.�7�z��
�G�g����i�u���G�LZĞw��mx�������j�����F���.U�N���*&c�������j�Mt�33A�+(��'n�NSS�Z�4���ף��Y1����W�V����g��BZ�R�*�S��̘��MFL�Bb���ɬ�[�A����:�M�_`�0��з,���<���nblo�\���?g����˗k�4�svn�ݙoiwj��C_����n����WPP�3Z��;����lM��DvA|��	�x���P�w��8�ܚ�d��4��j�L�Aal8��;i+kk���k��ƀ]q�<�p�z��9~nQ
Ӛ]^^�.�R׼	��}�	���2WCK�s{�����!��b�LU����܍��)4���]d�ѡP㾚~�\����!5�Y9�0���R�}X�щQ�$�\tG/V����\y�b�n��/$�����*���(e[T5:j`ii���a
L���#B���@ 0{�=�Ç�>�4

�033�s��?���`�c���I����-���|���>bf����
�8,E�W彼XA��J�ttt��ř55�'҄��^�N�����H)�@�( 8��A�������O��`K��K~4�ֻJޖ�L�{ssӒ!��%/&.nю�澾>��Ztqf~�=`w�U�4���-ml�1�XTr�GFF����R�l^8l�l��t�s����dc�T�,m�6x Hb�$���40�~���Q��p.�E�[_o�������t�y2�6���A^_?:��q���"R�@�]Ee���8|�s@k���gΜ�,,Tq��|biy�
]�8��,%e����R�0�ǏǅU�q�.U&!���r�=�Z�V��זʐ� �`���f���y
Vbs�w4[����=_��{D�5�n��eddܡ�⾛�lkk�Y�Afy����8�׎��No\��]�
�-���ǘ��+ٶij/ɹ ���#�,3}.F.��I}x�wl�qNy�B��N���T|�^'��{{z�'��Gk�댊���'���M�ֆ����?�6���� ��w��N��qQf�S�y@^gΞ����U�����j=PW��D�kj�bQn�VVV��W�$r�\��#��U��M���� �u�1_H���Q�u�,���r���6�)��������V��x��첲�����}ǟ�0���%�	B �7��㕿SR~��"��X��t`�8�k�@�����U�CCC�1�S.m{K�`�/:�0nK^B��؁Ϛ���)(�0���ٖz�� t��8�B��7�J8Y��ںChĞ҃��~��w��p�]7�fn<��qs�\���o�?���yu�+U���y��M����_}4O{�}2PC;��=�}O)�7W�'� ���PTD���A��]c��Q\9��H���}#e��¶'�+A�|u�3�!�fg��.R���E���{��bAu��������� �2��U$MANE�����jZZ�=��� �k}�0 �
�i�Լ֣rOD�0[e�30��x��?2r�;N	ܻ�A��+��Q�?n/O��v�ݡ�CU�.$2��/O�-{���Q���.X���d��!@%����5Y̥
����hM��?Y،�or�i�l[�.!�dC�\Hs$��-I`yUբs�ξ�S�2S�����	������+�0�̫`�7��������}�>���-����7�b�e~���]W'�(�!~��%5cc���
5��`� L��}E�� �*j���v���eA�'''�nl�g8���>?±�ۘ$������
��]S]�h�WL,q	v�]V�]���h�&���Hxm��^
o���UW���PY)h���cr2=J����|gG=|�����<�*�Ȟ�z��p�_#0V�;m-SO����T�W��fF*���s]� я��ǰ����R��h~y!r6zdD����%�k#�U��Ouut�Kbg����;w� 1���)+7WAi@��4Zq�����72A ��f��e��쀮����06�LO���	��ny���0^�U�G����ʿTU��Ӿb����{� l3��f��6�5��	}�]Uj��`�Ż�����q��/�����ۺ��.^A��~e0��>��������w��L P�j2#��PM��H�� ˄:=1]TQ�i����w\�V��E�,�r`�Ƹ�T�"t8�˹��˝fU����r�C�	�(�摏�IL��+�~��]&S���q�h&��$�؈�>x뻑�����5K�jr����lr��Ν; �M/䕺,jem�PS�]����yo��UyS��H�}y�S� �똞�,%z˱���Y\|����nA �e K�Z��Pl�-=1��hhfFk���߾�P�㞷3m�%iˡh���~�6%}��������uϒl������ɂ|*�PB�\�����aj���{�0Z����U��; \��M�?����,�'�5���ђH��SƼ��cN��b3(D|g���Ǎk�	%VTU�����H,���K<9���ۖ�R[���YJ��#�C[f��b��?�}#|��9�Mxx � ��E�U��\�_%�~*9ۇ䂾�	�9�Z}��9ܓ�A8JG;o��[��C�4���3�I�����w� @�Z����C��B_Z+K�sj1�"����Y�@���	$�r�*uqu��fk�W�r)���XPU�k�K����"V$$�	_�?ت2�W��y�V<�����?�޽{��45Y�+m"��-�\�ِ���=~,����i�Ե����0�#��Ƅ���_eW_��OT6��ݱ='�L�������n-V*��!AG�I�&��5��U�O� �B'D���G���aX�$|�fm���������0g@@@��O�z�F��e>\�>Q���6��+ �2u��󞘘�}��l`�k��M3�
JJ!𑮮�Ԅ$_�	C��+~���@g~�8�.��:��&��Ę}��@�v�l��	��)R����=���^?�WSSK�:  g�^�=]C �K����s7XϹd��ɰ���I�.N..�N7��7n0~w؆/����~�^^�I�=y"�{���B-Vr+�?'�0�|K%ءH<���b/=[��T�A7��z��������zXsY�J6t8�+v47�U����s0�{��+9 cǠ�Y�ǡ��䯖.l
޼y��1U���dr^�\�tl? ��U�'$$ĠN�����(�eɶ�Zn�]�,������P�s�]j �(;��aj�Ŭd!X����>o�=�!zk���l��	����1�hLt�₾��[ �U.0�D*��/a��Q]���b���ѳ2F�*���i����r`��d�M�KJ��D\:&��e�)؊�S'R��0�f@�t�z�
����r߿��i�jت(�P��1��[����"�G%o?�����4�p��M�W>>>֯ƣ,&��]\\,�/�
��{z�Ԥ'.-?y��=@*�M�EB���O1��-<�,�`�svqwtV�mwk�Ӛ#LK��U��aX�&�|RZ
"���\Hhd8������C9�C@'��nB��Kͻ(�*�B� }��a0��Ȯ�(8��i��$	/WLx���x�k�}


3�{��{{޶��i����m&�i`�P�!�Zsps�-R}��h�GJ�C�=���9Nr���UE:�L��%}�s�#)�>����D� Y��+���"S�LnTcے��T����O:� 3r��Ŷ�\�I�������5�Yo�_;J`��u����&&�wk.#\�Ν �/�=~A51����Y��SSSS^>��w����J�����Yv�F������$%����Έ�j�X"쵢DKg�C퓯��צ�$3?~(�[���	ܼ�V᫢6�g[r�Q[�z���7ɫ)Xq�(,?ː��K��<e�}��KY9��EW36_�n���n`�h~����9Uޱ�L��ɇ�z@c˕#�++q�ui�-��un�J�a&�������YJq�%��<�Y�v�Ω��&���b�S�l�[}�%��9� tb�D%��Zu���ZὙg|)�Y�;�Ҡ��Gi<N��q=/m�C�^�j���%o1��h��av�ª2�U�H{�'a�������0u���h�\_ggg9`4�´c?'̾U��s�	拻����2���L��X�s=O4�>����X��54ڟ����h$I�EQ%I�
33se`Q�ϗ<C���#���`jJ���p�\	rrr��m W�u�>��sB`z��3��XG|@���||�SSS``W
KO\ aHHLNsB%G]O_��?�m��N�v��5kna�W�������b�qϿ/J2귘^�p���vR�
����ޙ��!0v4���w�m�Д��3YqFQr�c���>(BߨG?� �p*��g�V&��0��Z�H[���}�B ^�ms�]]\��S����	�=�7D�Z���)^l�2HN���O��!�MLH�*1�\z~��)���*j��B[�-o�'$iX���)h�|W���wYS|����#N1x�;6x��*:ԃ>G�j�!)(�z��<���Nj��X3��{3� h:�fv�3@o�����ڲ��fX��౅E���_ �e��x`�E%&�ْ<.�*)��p[n]�B�f��實���'%�Z��ky;���S����.�j�O��
\t��[���eg�:2�n R�v�@���up�Z��㮑���]�2�+-�3ч������V�q���w��sj1���O<�����������KK�jB��11����#@M��?�T����*1|�������ʈPx3������r�I����,љO8
��;V�ŕ�L�}���������L�1$;�r���^*Bu��%BG��o1�d�˧.IHH8��゛�\��<�[�*�:�s�f
�[1P�X�����1�T˼��h ��F��lkkk� �ް�~`�����[ECTT�Z 4� ��c���!w�0m��+���Gt�C#e�,��
�Ա��S�w/MzM��&;����5�xIsR VA�^�y��w͐5߰�a�JI{��0H��r��D��5��y�+
��3
�w0�G�M��ﻮ�����׭�~zX@�aDa!�R��d�g��\�A��{|��ѕ�}Bbu]]�.;�D�U�v���eb��ŀv�b9�����|�U�y��KL���rM��ҕ1�<��Q������ c�"���P�3R�����l$E�����!����}Vk�o����2����� �	�͙3g��@p��ac��^.$0�Oߋ�����Wϟn���S�'g��m�h�KU�8*p]��B�����e~$��+���1�v��6�T�^����z�~�U���d�����e��-�Ȃd��^a�T�G�	�u�����U:��$�S�S�����f�� �zx� ����A䶷$ �j���N����Z�!|�΁<m�7E�+W�J���*��#ߦ�2������Ѯ���V���p"t����h���
��P�L�3�0C���E8TQ(#/e�zJ�444D��O1�ʜ��|�E4N�ޕq]���C�ll�������AZb�8v�z\�ɩ�������<-�_P�n���U,E�lL'���Kt�X#TPX[s���ͥ_�9�bQSSSu�
�'%ţ���+!��|_XL,q�D�h�7 55~�p�Y����3�!G�a���yN�2��͐uQ�c�t N�R�]W #JKKi���^ +���;�XIp+>%���딤�kTa֌�O��{k�!�*4��4r��V���|�$"Y�M�{�Q�>pK��f�i�gYYT�onnv��eA7�$؍�׊�/ʎ��v���4KEz�{���qm�#������B�.ͣf�+���j6S�`���dq5��rM�}65=&��8��]йg��� sVVV�>^���RR�@i�]�H�������6�6@� ���Tn'
��HCڥ�
]�Zzz�6�����g>��:�r´��o��\���$L�;8�
Unzk���94�hG$S�_~u��R�Y���B�	��3g�f*DMMm���>����%���ٙ���&X��4��� L�l������`nаj��WD����[:���'h��)  � ��0�=?H�] ɚ!S$J���-�&A�+]㉞��1���zz�LF����ssOd�����N�����aX�)|��Q�R���8ѼM0���p:���߿����*�he�ON��@���e����Yd�QIfay96��c����+������⫝̸�[w��JU��� K��]��0(�����yYZ*�z��FD�ͭj��Z^[;n�֨ԥ�(]�)�'��I-��4:FSl��ƭ[��+* �}�}���(��A���6ff�<������8�l4�5K+�(@�������b�tu��"���fdRu<��q�~{�q���/a���}�@(��|���q��6�x9ɃmS��}�ОE���_#����pj���c� j�s�Cs���!fj
ΖZ����7����F ��4/h���&�Aj����M���1芶�1��]�0����r������r�LP�T�?q�/L{cc1*7�/X�����}�k^�6=P��H�vv���z�ͭ�b+:F_�sEEE�O����=��&<�z��mv]@|�j�[�����	,� ��(�J�o0����m**� �cee�	�6���[�@��l�k�0yfq@����S��E�KҶ6/^�(/'���,,����/��8ඇ�K�Q�"Ҋ'���΢3�lTe���z����	�w�ϏnBEV-�Yu}������lp}��ff2
\�\�_��F���=}��Lןm��f�f*��v��%/k����SՅ���ܹ��eK��}�穧TttІ���x�<���l��Fl�.1))ڵ!������R��]����U�o��S,PNCL8���^�l���BSӒV"C-*�ߝ/q�%�$*&V��4�krM�!"�`K�[2�DmD���4*"1�������2KZ��$��S��R/��Δԁ��t���#/&���6��֑]���ԛ�I�����G;���ε;�!=.�H�0֏�3%%�sE%�Y�KZG~ˡm�v9b4jw�*��k�򼋸�I��xf�ًE�
���C��[p8��5������dn�j�g��n4�ޤ����Ɩѷ�O+ۊ�T�66�|�kn1U�i� ���̆Psbb�f��d!-�����FΪQ��n���&%�ky	(++�}�C�C;�Z����pBJ���?��u�	��9�eqs����ƀ�f�1�h4@[�e����_�<wFPP(+}��b���UY����:��iFG�m�=y���e��>ꞺK7��\`�}�^� G$y�./M�\���9%����a9��_�!�J3ӳJ̾VX�����,�T�o�����	(�
�����Orm�7��F|�@�Y3������Դ�d�E=��ɋ:K�ϼ�\yQN�{gz�V�RM���c﯑;�	Ӯ��C:��<H���cS�،�;�OLH:��kT������co�MW��}��;���O<L�ju�&�@~R��1��/(�E���j�$�p@`�L��y�+�RQS�i�ο�U����G�F�M����j��w�Ѓ�/z���SZ��ؾ�]� 6"P��L�%�-L^���`ұ�����*��˓hdb>��M/�XG
�@��4�g��	g������0 �ޝ�$�Yn�{��QE��:'���]�0k��"��G�3�7���!� %߹�������fC���!|�.1��_4�[FW-ڱ�ۑVW���G2������@E"���q�H��
t>z��y�z�j;� �1��t.@�$�һq�Y��
�X�\�P��ΝE7p�~���V���9p���p$Ͷԓ��R�NI��oP����������j@���~����f��ʙ�4��Н��5N938�x�ݥ�2�+Q�X�=\� O���e����R��������%@�!u�~'���钘�?\�U	h���_��y%��m\�ЩQ��x��w���8��2z�o�pl%����3e�+�c����@��5������i��C��Bf��I�U�M1�w�(C`[О��^���#��� �[��WW��?e����l��A��d!:������Q�[ ��O5�,.�\u��^�2��!��EJJk���)������?�5��옧��J�@8\�N�(E8���Ã}�����/� 	%�-%��VSp���#H��[o���7'���ɪ���õw�����|s���+螺��E�!㯼1U��!�e��Sb�!̻(y&e�0/&!uM �)�g��Ɍ��99rPl�_��u���3/���;�	ͽ��j�xG�&�Up݃�S|||�����@iD	T�	�E�,}��="��W���2�`��� +kk��h����j����$q5H]�x�V�#������9	m���;"%p6�SE����洀SvZ��4���y��mX��yԖ}5�Z���H�;ą�%w_Z6��&º��氎�yɏ�Ǡ��Rgi}��8c��X��ǚL�w�l�������]�	�?��O���ݻ��y���>���ө� `����6�u�����PV��o{	�}�r?�����~�"~���P����AQ���p�b����o�n�V�9@?�@|�L
9��4���0=�1 HCУ��hU����`����T���� �������ڑ5l����~�<Q�N���b�����S,�7�f ~�	�{:�Q	�-eδ�>v���](𨥠,�����HpJ�t��~�����F�ƎN�������ɗ/_�P�"�������$;�+�\�����MRVp�]��|9"(��v�	�hL��)�i 	+f\����4����J�����^
��!l�.6z='��!�/�2��RsXr��Y>���u�(�������ͫed�����XJ"VT�;9�~.Y:+2��V>V�y#�/LSej��������-BK�)J��o�^l�	B�kXX�TJC옗<�rr殮Z
���'yCQ���Hڅw���e2x�0n�5�j6��#w�qs?"aT n� X�h̦op��u��2g=0T~ڢR�j�ͅ�י�^P���^[��_���7�#.>6��!�w�Ssc�f9X�'u=Ch�W�-�F��%�`�i�>k��\��^���b0!�,X���"��G|������3��6�B����Bծ���ܸ��%F�ܼ��zQ�x����'̀� r3p��>�ٹ�}�j��2�y��HB���>�ɘ��h�aȘL��
p�P72��Tx���a__#kR�t��{Ν��(m__���w��i/n_	��X�~��D:�  T��@���bfy9���"����n���W���T����fؤv��/[�ġ����b0�N߯<<q��j Z=P�/�����jt�9�|�9�`�Q������q�@�i���q���7�
s�\u�3����	ܒ��$�ٳgK�u�7���f��Mjy�h���Z�z{�W�c�lP�}ea�WK��-:��(���75ͨĐ>d<86fT��4����c�x���t�#�����*��T&$y��L��l����/��D�d��B
�ۑ�6�
���Ϟ�rkr�m��b�ihk+��?0`�`H����3L����DB/��0]#���"1�jQE��;����Z� �=wj������S��f8j�����2��M�=�B�N�s��yG�8���d��5�)�琭��~O�>�U��p@I����� j?-���-Oqz15dVIII��d�������
%E%%�*�j�#y)��L���WAr�"fps�[0�R�d��Ah;]ۣD ]��Ȝ�Bද^�������;��B5#�C���44�(,�@@�=���p��)��>�[�� ��Kl&>���������ǎ�	�;99���9M�l��������R�E���]�� ����@ ��YY��W/���>d2zhn9'}�0�F�����s).&&F��Z��]��xC>I���[T ��iu~���>�	|��]p�9bt� 2W���q������"۳���J-@���� J}�ޝ1��'��B`� {}�'o��V-��$GL�}����ӣ� �p���	*�����oU��9�z�n�R�PھrZM�*Y$���se���::���J5��B*;"MMM������חڏK�T�����N�����|fer�,>!A�ȍE�m�	���_� <���?u���W�\��,G�4m��.l��[�m]%�mj��H�B� ��6�U��V�S���:��x����.��\h�@�_�H��m`;U~�U/��=�~ku�K!-�^�)Qz��Rmڍ�4Ad,�I�_���^]}�R��OOVMx��dK�#vT����1>+"Y�,��Hr...P�M�Vpi)�5��(�=���1`e[���'����)T{���A͏ ���aյ�XUr���P��)�b��7��!��0E���x\85H�&e_td(�^]�uWv��e����^_LVV���˞�M����[�ku�������&���)�sձ��$}#�q2��nͮ7�oÕ�(�^v�1Dw�P�s6�^���ia�[�������C���ܓ�O������߭odG��y.���4���Y֛�`o�n�)D�S �����wR�ڑ�ua[O��<����]�|ӁR{iP;Pj���D�c�GQ{?0����Ϫ<�~2�T��9%��ڛ�(]�x_��bh[ڜ�g��z��췧�E���QQYy=/�=H_���G`c�<��3����s�}�X�B��f�N��Tt<u�8}=��� �b��� Mkrrqu�b�ff����4.�J��n�|���;; Fk�n\�O4�hU�J��BJ��|�YJn��DeT��V߂��9'��fq��ZdT}������j)��Ը�m��� N���EE�!��2�)à~|����T��ږ�24b�WI�� �O��>(��5���IE��*��n- K5��1�2������f���X���nAZ�����(͟�`	�t��x]�g��v[\���Y���z����-",H��0c=��\���f��o����/��B#�H�|�±���\$P��&�so1ө��������ﾭ�8�?V��G�������gU47?���>�"$�~���eSk��/�E�:#�������Ǎ*��O����/,����.�cw'�������������-�?�Zш}� O�^)ԯ�;����W�k���U�G%o�~���֝��b /q6[sWd˲�yxG,�8u+��i�Ն�"LJگ�|���Vn�JBA��JGR��g|��܃�O��0rg�!�#]_[�Y�!#�����dmnn^�*����,e��,�����������ϑ�XŻ�9���e�`UY)h���P�9�3.�ff�_�;?d;��\�K���B�J��z�,�}���"���tbb�ז����;�Fcw1+�9�c��h�l0���(=�l+�R�6~e��X��{%�����/sx)+��(����"\�'a���ƾ�p_�;�����W���	-�4����8f��Z���Ƹ�����C�~�@���moW�;��sg6ҒN�c���:�s��\�1)���	�Cfc����S05Uh��P���j�Գ�¯<��ا� 4N�����ڔ����w��U�������棶�JT$z��HUe%�>���\�6����%�4e���NB�6�؀�II�h<�B��@�A]����
/^~��'��ٮa} �h\�����&�P��D i
$��(�D�4G�hS�ή0J�&��J`��~H:�pw��J�rf��8�*�>�'��,*��@舏���s�xd<�0Ω)����+Uq�WMӽ�ܪ89��H#�9�?Y���>-,X�e�M�L���*YP�����Ynh�0�c�u@�h�d�+UϚ����0���� ��m�A�Y�U��"g���o�%~�BA�K��������D��tus3W��X\��O�Ki�Y,PU��%j׷�����ӎ�K*���I��(ی�T�Ͷ�lo��4K���~�=�K�?��*���c� �DB%E�T����n�VQ%�K�^@:E�DriP��EZ�����y�#,�����w�̴��0���$.��|֮l;ځ���e�����Ǽ�ԏ�+҂��u=��g���:/�;�(�t�Q_0���R���z���ME��mCCq���i��<�����E���I���E����ʊ�ү���׸�Y�o|Yܰ�C)��]��6OO{�p�<���tՁr	��<���F����Ys�����<@�B~e��c�*��0P����h��~�<��_�1"v��uD���il���2�����q�F������j�8T�-ܾVXV��h��Rs>�Gk���̔Q��t��0/G�iO�vs������,l�И�ѡ�Osm�Q6�c� O�
�눛�؟�#�a�m+9���׹�=��Y[Z�P��ȅTtZ���{��]�I'((�m������S�����,��$�m�CBg��uH1��o���`�ײj�{�۩`�r�Z�e�6���ܔo���f�|��2ѷ;jjj�s)��N����=*O\Ěz�����\�`:z" (�]g�P���׀Ic�/����g�]���=��-���
eܹ����:���V��K1���oG�"Z	�0GGjD���2M�B��oD\f��H}�b���P�̻�Ys�����q'���\/��Xn���n�W�_WB�������	'�bEa����}�rR���a������0m��3Rs���o��X��p?�G3�p�Up �++�ş�M�[���[1-�a?��,����������������P>q���2���P�&��95sE�x`K�j?�����ُ������emm1��>M���MD�����b|
�-��]��w#�Ε�t|�,</���<����U);�|V�y�f�� ����e��.[�h)HT�RGlc�9ؕcaL!��"<�UT8��=#-��NqwBL�l�o#�0:ha��t�f�x����l(�DȖ�*�3�����Wfg_I>�?v������U6)IzSܶJ���	^�:s��������h�L'�ώ}�����j��b�<��zl�n��R<�3��Ɣ��t��S��jQ���sL�@��3��՟���W|BMI)x~�֠)��-�?v����ʬ0�)A�0�&r������I���1.i���������sN��t]�8����K�!c�[��#���6��e�r��&������3ĝO6vvJp��~��[��b�3o�v�
���j�툅�AYy��l����8�Khy���t����{�V��ƞ������;����x[SSHIIɻ���(*�͒���=�)�9W���	�sFje�cq�c�L�&P]��3?��6/t�8=
O��ģ&�I�<��ׇ�����_��o{+�PKv�a�R$��%@Q-I�{���6������]�T��u�����,I�s�5�c���e�Ԥ�B#�N�[&e+r����~�8cL��cbo���mo�;���������Q�zŮ�ŝ��HM�2v�
I04r�W#:Ú�L<=u����a�����qN:�喕E��;����Z���C{j/c,��o�TW���r�}����7��K���W<��I�6u62��646N.��F\�ț�!�ݣ�Ө�L��(��ɋ!
/|T�<��U<�ozq��a<�cXR[ו�can��2�=ˈw��|���4*��5~	hd�9��L5�i�ݯ�A�"�B5�.�����^��.Pbn4-m�^u�|�,y��!+��v���C�eZ���&Oڽ���=������x�G����{%v���v���\6�"��~����_��n����)�<F�*�c�f�Ӕ�yo�g_Cn!���wY�gM��������z�Ь���c9��`fz��X�8���2)<�X����Ai�K_H,���T��	�(�5��m�����>�-�E[LA��ED�a.�� �muH�����l��&x�̺��	
C��������j�\U��c���bt�C��R���n>B� ��W�\Q)�@7�)���^�ݜ7�]�	�6v	�f�X���T���*Z^v@N�x�<�cÆ#���t��e��X��r���U6���3֜R����'����S4��M��]Q�\	w�vI�V�wЍ��q��I[q�%�~B�jr���7�]K��1������=����f�jg�B"#Qw|r����͐�/��s��,���m���g������힒���9��F���h�Ξ�Ԫu	
�w�T�N@ԁ��[d/�/luF��ߛ4�c?3`�l�������Gd&qo�c��n��Z*+l߀aQ���i#��^�����We��,[�����z@���7&���fA�ɱ{+���
ov����J�W���\�&���pOQ��?���n��Y�i�R���D��a)�5�(�� ���ی�R��ʴ���=VV�ޣc*�A3r.���G=ϓ����t���9A�?5V�[r�i  Ԛ��AbĀ�+�dd�eƛ�8l,�bDʪ:8(#�ݭ�ey�Ihm��>#�Բ2M|�G��RY	F')�^4+��Q��.��2�J�&�z�Wh7�����c'����z�ڿ�b4��-�G��6o,���(sjk�QB۶�1�I�� #e�V��t�xe�o+rv����./-�R����sv{J���`��;Qc�R.��*��,4���(툞��<ԙ-F��\�X��"5����8����@��|�k�`�#���F�yu���δ8f�=;33$-��#lz�7d��l��vw&��MuIRLaC}{����ΎuD���0���g?M���|�i�������������QN�Zݨ\��ܯ�,��5"�(�֋�&�Y<^�У���	)������xٹ�4������'/l�c������Sl'�i��yrr�y�q�����¢"T�6555vw��>w3����?�;��U�������w��1��ev�@��<�zZ�i@``r�5A�/���m�c�u��}QTZj�o�l�
�H�P�P�h�����Xf�g��R�����}7f�3�eb4��{���L��o�C�,e�A�x�0G5}�]g�C�?ߞ��E,�q�x�۔[D$��D��F��\���=u���v�"��;ZN������4���K>5�G{�b������o�����2\镾=�����e��(t�Ǽ�w7Z�\����͛f�A��5��n������̏�X3�<~c}WC#RUU�Q����-�lx;�U��\j=�\���8����r2�v'�����8�Oz���Z^�O��۪Z�+߰���~�䛺���������*��+��	F��E�5��>͜u�[f�)&����@��RQ����QS^i��d�5O��|TYQ�񝁴���c�_��;���	��ѳ��U�dj�VXX���������L�ի<zs��"#�
8?𽩣O�<�ߚ������-��̗����"�	&5�� ;�73K�2ibb����,�R�f`�({����[��Cp�U���"�!��TSm�齽�t�.��d�ȤYx�F}����Bu��I�C�n��*)a�ïNb���[�s ]f`N&�4����2q���p\ ?c�T�r�f�eq$��[���")�Zͼw�5sAqE������wb��L��l�3��k�Ȯ�n�;/��0l8�8�me�|��R�\(����$$$>[?�� �BF�'Z�to�����x��QK�ַ$l*�������$>~6��ӓ���S$/����A����dWx�V ���W�M;}����?��j�UL:� O��x_��V��&U��$TuJmzwG��~�����Q$	j�t����c���~B�Ǵ������e���]�
�G�.=��}y�r
:�揉pp����KI*�T�o�ʜ��}tXZ�K
ڦ���Z�Ś�<z�?�؏ .���=
�����CJXl=��5��� 
A�m[��A�2�622�ŉ�皂�\D��B��-,,xʮk���O�u�U�]mX����9V��)#�VH�1�ɡU�e�g{��a7$�g�͈��Eaa�0V���0�y��gϢ�ͳU�ɇ��s���9M|�'^ԃ�	���sC��q��{�W��>O�D���$K1xu/m�������(x��w��f�.�������5W�ޭ�q�bHF�и�J����r��ױ���؝]\b�ڗ��8�����[�>wt�N�!A淉�q����UnC7
�-�Vg�@R��]n��	�7����,��]b<��HUY9)Y*�"FX�/O�k'��A������d�zcD�Q����u���ǜ`�RIW��ݯISJ��x-X���s�˩�����U��	����Լ�ٱN#��o���Z��mm�W�ၔU�X3��h\b;�_ �U��Q�M$�9ݓP�?)i'�^�}���f/����ZL�]�b`о}pl��C�`����Ȍ�!q{�z0�}��i-��j�f�)�Ú�����W�c�2AS�y$2�'g�/2��X�v5g4+;}I*��Z���zÞ���	pp�q�Lp�69 �د�%s�7��}m��R�د��Ƶ@[����m�Ģ�|�śqk#Un[ŷ�w�#k�Kk�8�44,[�8�W\�ml� 1VA6Ϡ��\�@�x���uT<��F�d�T�}����q>|>.Zd;*��p9�_
SiX�|4��+�s�SANw��$�ߟ]X(v�J�+Ӊ�Va& �WUS+�g+mw{�'Y��0�s�I��v��hK0������=�ꑈ�Z�'1��Ͳa�] >�p�@��Դ��o<5ϞnK]�e�Ы��C��������r5Z�d����U/�#��;�_]��kkޑtW��H���Zts"lko��s��#�\�O՟+��;G?�,L6��%*�Dp8�4�-���ZXY91�<>�m��f�l�e[,�қ�����.?���x2\�j�K	**���.n��Z4D�/I>���t����im�<U}}���!閣E��k�0��7j��e	��=��-y��*7�y"l_����Tk�$QF�%E������&�����@�mO1�j��~q$eF~�i:�+�㑸܍�_6�J�D0������<FO��'�CL�z�hA��&�.������:z��"g�����L��c�Tk�Q)cj��1�2
r2<�[�3�����W�K��z4�Hݤ��4p)3�@�Տ���i{�ؒX\O���sa�u�7TOO��j˛���1P�,7;�;U�������1����`$&b?��S����ۮM�)^��yRE\�˪���ޭ[Og�	��ώ-]�Q��4V�kg���-(�kje�ǲ�jc�~���A�X�@�Hq��u��c��xC��#�ZK�єR@pW����,i�6N|�~q��Ѧ�@��o�Я_�����DyVC3��ں��`.��6����u�����3����?랇ř�~P���4���X7�4����no�'k�����@˯��	s���S���Y�߾��;L*�Gfe{_��r^�c�;�=(�G��R�����;�o�&�T�]��>M<�O�$tn(�(eZ�3�*6Ĩ�1r��m�tt�?�1ou�	ƋyH�8;�iRs~>�-g�)�Q~�/>� *&$���>k�dfN+�>!��Ͳ,�}��>jٸAhٙ"�74��XD��%�7O��JBE����?к��⛫�����K�+��r劣��Hc�^>*�X[[��cRCM�B҈ʳ���/h�dxʤ.�<�Y!���o���kh�"�]$�����朡�TȺ!A��+��k��Wk�c�K�K�+T`c3�掝8�eg1}��4 d��Y���(]��g=`l<�9߰��Q�E�cH��!���gu��Ĭ��W��ӱ��� ���R����ɒ����><h�x��\'Z�0T�N�Pi�K���܍!��Y55#�G�?���s�JxB�|,���eH��38�G'���v�߿�TB���G��k~U<:�|��kۥe���JГ��7���)��Go;ma��֭}re��}�븘��լ�ޛ��a����&d��y����ï���B&�nS)�����:���EO��������q�ؓ�:ુC�Qge���*EŪX�5�T���0���0A�O,�m�zp�p�YK1T,�=
9ޫ�EҠ��C�v���+��%a�1�<nl݇DjHK�2���lH�fw���[\Ă�0��kؗ�#�����,m&7�7b�I�V�Z��K�7��]�qV�JQ�>5��{��A����V�HkZ�~�s����Ou[�06|�MXH���{��_��OMx�y�!�	q�dA���7٥��n^�w1QW�P/k�'**ʧz��.����"))��;T�Q"����v��Am�t�őj���Y���*�p
^�޲�{��o�L7�I�#�2EA���[`�����J���KWv����(y������\h�`�T/�b��N�~q%���S\z��O�����@��O|���m6b�$W&u��"����]L�A"�=btG9�E�d �.��"������M�?�U p�#_���^�ܜ��fH�k�C'HHt=f�d@�Y;I,����@�^�:��5�`t{�֠]|��`�XM_?/R�]����۳337"����V��;o�@�ϓ�[���f0G��;�V2��w�n:N����f9H�]��{b2�6������&�$�<~0;$$�N�A�������#qj�
v�v�+�����r��au�������7�YV��Y����]b=�������z?��^m�n�
;ם}�8r�H��'�?�b]̌�V�5���ɏ��W����4Ќ�1�b@�6:��	κ]|�c��cߣ�2��,,��H*�izT]]�V.w���E����[�,�����n>\�&W���H�Dc��Cρ�E��oċ����q�� ����bȫ�"��%��>��&�7��ïh8A������<�$�����a��MO���M�����<�����ih#�bUJ�6؛4����:��Br7;ہ�,��a�r���	�~Y;55�O���%���ѿ��H��(��}{{!M�@��,�A���T�����uP����3W�*����������&�d��h~|R�5�ݠo��/��C�l�f��0|�=NШ��ᝋ��mlwZy_sZ���*9P1� -ւ��n
cu^�u���d�G��r��ɒ��E�]<Fe��@.l�	�'w48��D��S����Tma�&&��MRQ�Rg�XZπ�!�%��ǄYʶw������
~�ȡ�(ݶC��5d�|$��.D 6A�C>���@�M_��6h#P�&L�UUC�T�C�w��E�x���'!���u��q���ֆ� ���{hh^���)e9�7����}}
�|2�,�	R@@}[ܨT� �y�h$>��5����	H9��
�����-LHDDZh(%mv��#D�e�g��:"oW{ �վQ����O���近G >�n�S;L��ch���*��wP�2�@�G(DT�
䀋�t11I-�*3v"��>�`�ӧ'!����f�� j��s5���2�O�Y��u=S������h5z��>�����P�;MA]����
?EM��{�3B)3Z̫�J�ȈϾL���_Q��?�&8��.
vJL�e�K�G��^��=�I=�k�n�KUK�	�q�5�WX:oZhx�1�U�,x�sy�E!��׶.%�e�����0�6-�$/���6��P�A	�����v�4t�A_�a�*��ش2��Q���ª��$��A���õ*��C�|j�ddd����ՍH�/�?�;�ޭ�aa�F�����U����0�/�lԵ#�~���v/�8W�Sz���� y{LV��(����	H?JYII��ʠ���mۚ��
g\�qY���n�]kq�G�!F�>�f;w3�qP�F�c�b|(P�-�RE����B(�]5zA}��'�ugy�L��a�j��#7=c�m�WV"E�-8=��V?�����&�7T
�Q��ܒW=���a6����ȩ�+%�鑜���Ⲳ�bx���No��s�l��B1V��h�?���׳k�׽���^�07b=�\���kH12��&�u��c�W2]��-�w�dK�ï$R�`�#��a|D�,y�l��z���"//���s�S�.���Iru ��?�M%P����f~��-�����)2j$������^,lOg���r�"��a���03q���F�XP�ϩ���g�48=���޶�jl��U�g���H�@!�ǯG���:g���&�O{M^1�7^�����,dV|�U���BV�3N�m1��:���u}U{��d�+y�U}���^]3�:�pf�KBW���M�2�s����]]F(�*O�:�QT�l�u �Q	u��M��0(6�`�^�mOM�"��C_D���A*��U��y��щ{���7��]Lk�I�9S$uPpw�W)>��N�;�<c�݋��]J �H�'�9������ˠ�+#g۹�)P홊�2��z�y�%�A#M�BMk���xC�����\O�b���c�l������p�����L�kG^y��㋰Ʈ�4n�z��EL>�t,) �$�]���m�����^$�R��H�wyⱢ��V+y㧲6gI	���6��ߗ��~�ZR��s�q��2��<B���o��D�5ۭjD9������R�ȟ1���e�Cm@D&��]���Ў-��1<��{��}�,2|���3������D�)XG��]b��ø�����F�62߿�T��F��O�����􅪅�/u���l*1�E�(:��K$8����N47����)�v�{���n��'��뮫՘�El�I�y�%��(���Y��Rq6��<޵H�G�,����-�������1��!i��O���}Çl@�j�C���|�}���rG��)�,�2���ÆdbfS��9�];�&'S��P���R���ģ��TT}��&�U����׮�,����uE=G:�-9� ���
R�k:%�3�ttt%9�K�uw�;��kG���W[T���(����*�+���MϮ1�ʜ��-����҇{�¯2��\������ȃżC����| �O�&��D�	�$}=�sC(d7n���e?DЇN�^�j��#$��hx�
�kgs������̇��-�̎C���l�!���3.i������>F�%���Z�׿��3����ѕ]�xz3��C% ��DSXޤ����^	�R¼lo��x��D���ɳKJ�Q�XG�1�VR���4X�Z\cjzz�CRO�G������v���-�֎� �|��qJ�QWa6�=�������4���X���Ħ�_�V��q+�E��k��,Iz�))a�ԲfģKWد]�Ӗ���ةspo�&lo���r���������&rYN�ѦD�������ؓb ]4⦦vW��f�Nw���|_ܐ���!�&/�A���!��K��g\ބ����k���$!�)�J|�T@ts`|)$v)S(�A�.d��EN5��Nj"�נ�D��P���[?�A��P�8n_D���ϣy�X�<�j�F~S�����=O���wuuѵkiq�Z�|�aucuH��9V���h�{�1Tink���ݦkg�r�r���&Ĕ��C����͇F�I	�;�虳�˩fo,l�ֽV�^��� �2�ځ�9ɪ���s�#�ϲ;�~Pn�B�ɉ����`��u(���w��"���0j ��}��X�W��Dy�����|�PXG�ȱ���y�f��r��t�x�|ޅ%.�y�ł�̘������bcem\Z��H���(t[1m�<��cO�:�sU,*,-�},�ש&�@F����ܷ4��&�X*���<t�آHgum�ajm�ڍC�����#��=��X�ϱ|��^]�R��iuK��s���cP�ib-�����z�pIN�U?W2٫J�e#�䂝�k��h����ڰG�ڦWf���wg������g����-�`��ܜ��wbna3j��{vi����ƶQB+ݛ���ވ�� r9l���������֦������'''�U+�
�bx[������d���/����H�����u�2����\����C�6�
���0;���a��e*��_����<�#"F���z�w�ė��S��c��SuDN)u��fo�p@>*..������Nlڞ�{�|����Ҏ���EJ���H}�!
��R����ɣ#�ns{��h��w���Ŷ2$��+�t����V��&��JF��9?�̮�<���87"��mP�yֽ-mmΫӯ�*��=*�g�'K
��
�Q����:*?A���c�_X��QR�|�3�Cg��ϟ�AS������3A�%ov\�qs��$������A����d�l�f"�J��s|����D�OsG�BD�.> �m(lf�������ܽ���cḿ)���N+쒃��[<u%P
%��̭�R�w�K��Z�Jm��$0���M%�=}i�1t��Z���δ86LI�F�m!�	(\[�Y��lJ�t���V�yΠ����sssׯ_o�X3k����R�ib<-�E-"�'���Ǌ�x����]�i�v����	���mݮt%���;X�*�b8��|U
�����Q/��LL�Ɨ���o���â+(ZW�H���(�|f�{r͠&�K��M���^���:퀇���%kO��T�ѱ�*>B'�$������bG:��eoNAfL]ff&gC{Eee�㴢��]\ ��_9���
��p��d�(,NMQ1�xX�#.�(��%� Uw����P�*�u����6��0��sӡ�Y ��<�q�*rz��o@��,��W�M}+�ڰh��i�Nގ��W�i���+��^�-����:�����,��G�Cyy�U������?��b<D�9jtm���<����&GЂ�m�A���_W=�
ʛ��De�m�ୁ���RI����$�����4-��݃��9K��ؼ����Z�S��כ��8Q���)s��R������2Qv�)Į���Y'��k�כ����.I���/ϚѫtQ�X��H<>�mmD��[j��������������E'M����Ɠ�.g�O�\.
z��Y�x��4K��M��o���:X펌跰2�V���Y�ۚ��@?�-s �zK��g��m��umD_{c��9\D���O���f���UT��0����3��׿�p���������6i�W�fR~2�p�KM�B�^��C�� ��7�kJ���޺�OCC�~�z�u5Ȍ���V#U���/f���tp��w⬿�>1��}�@�_�OC�ʅ�jzz�Wi?�Q�y���}~��i'��$x.7=��m�"��LNNnrc��������� v7ޕ�=��a�»������3P���u��ug���q��ܾ.�5^y�%��V}vK�������xY�ŗ@��Õإ@`�p������bܨh_�]�0!:��|��I޸�7��f��A����A�a�MwB��/ع����v=�)��7���Ϗ��.Z���N������Ac��7�e៿s��{w��o�-6=)��&A�ƈG�:/̔M���l�\eK7t�\��BK=:�9�ds�{�_�ԙ3s��������6�cbb�b~NMk��&�pŋ�N��{�J���Ǭ-�C)��<�+580�;J�g&9xU�?5V�о��͡�/���Y`@g:��L/���f��}_�+?�Wڥ2�J˪R�����7���9�[g��\��a*��ՏL�����2��yN��G[���̌�B�Eii~��� �y-ޙ~��YqFu������Ig�6�Ѿ� %�**6��R?����`�e���Օ�����8ѵn�s�6q�Ѿ�+����>����4��}Fz�|�J�^���ڭ�Ze�N�p�lW:����c�:��\��F�=t�}8�]�u�Y���.��׌�>7��[:R�:�/��.�������g�K{"�[{;vZ|�m�mt���E�����(����~��`���qVNě[bm߾�O�Uwc��	��{��b��!���,efff:�ΥA����v�曙���*Gwb�Bvx-{g�
�|kFƗ�zw���F:�u�������� �����NFG�%Q���NG� �n�{%v4��v���o�/���e�4���Օh�D�7��3Ef�3����H����݆{��rdm���4��4`s�A]=BVNn��������:�稩`$�ց.���TY�ݑ\[[�_��҆I�TIG��}���
��f��+]�q� ���N���LZ"��M,,-�F�=�}!�rn.V�,I�
���F����X�d�/�M,�b�{s���jG1��wcgc� G�J��g*��]O4��'�����XXh��EK,�}9ō���`�V{��xԠ��������bu"L�\�~��?:$���^|Nv�ΗHPLX��ߦ[�f����W=�����5��Y���5�)J�Y�M��l(��b��ǧ��Xl�B,�`����/���z-�g+�T�����|��[,Q	쬊�I�T{���F�"�R�->>�T����/���>�4���NIKcѫvW{z󦞞	�����̣)Mү_��U���7@1�ħ8��k��Ҧ������ u����VW3jk����{��$�?t$KY�G(%�ݠ�oő�ɋ"�zBd���NW>{vXt��Bl�aj|'���ay�e��YS��ٷ�� �%B��Z󝛛;<""0jݘ��퀺u���ׯU55����������9obV�^�a��f=
r�C/�x�ߴ�����n����sb<���w�c�SQ	.U�N�7�g�]G{��6���Lh���ӧ�l}�3p 1��.��c���;�!���#����뾻���N��<�YS��X������
��Pr:���N�K�jjj`&�y���;�n97����G�=e0���lll�� `��g~\����oacS��'0)5����(N#�p5W.����A�i<|�w�-AT-�2�	���E�/�=�fu�	x�9O� ����P�}t�R�F%��ƶ���l�6�[�eLl�3�K�	㭅�jKl���J�D-{�(9���������G��Ws������WI�gii�Xp.���P��GO�߹���'��Z]]�GL��^^^�:�
vJJ��6��d|��S:"E�y�h����SDѨ�:�.kn$O�:>x"bO�Ī#9X̂��V-I�b��h] 3�X�i��Y�%r�I�Kv��y3��ƦW|E\8u�b%8��.P����q�[[[��YA������_=��	!!�ͮ-롓\1���?�|A���ķ�<�}ţD��o��/����e��p�=00l�����Q�R�b����k���gFm3��#?/\%�&�,���N���]Ď��ُ7F�Sm�h{�.C!�Џ1�\;�����[���]%�#�HtvuNb{{�����e�d��[fc��t�����{IN�z�B-[�Ƨ�����
��}"D*�����3YEE�	�4�����=�t�C��� x�ut�TU'�K����e�'����WB7��9����:	�ekD�]&)ﶶ܏~����g	�!�i�C�F8T�h�í����yz%�h� �KԱamyQ������Tx(��[�n��qJ�����H���Q�!]!��'�d����ߊ���Q{Th���TZEgggx=GGԃmq����hy��tJ:6
f�aR�����#��9���btU��=9���k��X�'�K��Y�y�ή��g�Kٕ�:���|z����R+Ǯ4�L4�;�C�������?���>>���0U�$����CC9��.�%dXD�׿����N�P�vY+z��������'K@P%���
1w��2�`�8P֨�`i��������f0PVN�'��1���7�԰V�HhҞ(���U�ZM]}���R��XmvU�������g3lbj�b��W�§�փ|(�{Z�h�f��?晲Ā��=T>�u�dyסj���/d�]�_��B�paa!�꥘+>	���k�y�i�/�C� �f)����h�Az��2zKB�WgE[���T��;��(s���nO����]X�|��;�c���|�k�]��}�F�Z�&�ɩ�
͎����<Ro���m(�[3O$9��m�;#%�|�T'�]B=(vm���7Lk�Ck����/ c��n�]�|y�ZAʉ�@�/5��l�+� x�.Y��oU�n��|�v���Cem��� 7���42<d���Б���� o�EHp2���K�����@7��u��3�}{4��U5�Q�����)DW��
�'��]����ֹ���Y#�'�ۊG\+J��}J�d 
<��y��#<7n<`ڟh
������U��E�$��/���Z�?x0MO�K��	��^%&���j��d��ի���Jq+��o��{)&��nmo��C�	�@�G3��e�.��먲���h.B.�5>!�oD�t�0��q���7|w�HYeȫyG�{�ރ�^G��@�gٷ�����m����,_�j���&��
(�씔/7��������;M��ӴT�X1���^j���I�q��AQ�\�ڑGdK�d���v&�Y�29eH�߬˄�"�z�W'���h��8O/??n'q��"e�u�M�]��."WNx������|Ƅ4N3鹮���{����"��K(F�G]	�T��bh�sܢ��&����1�b$�(y�4������*t��|;�剥;�?ٰ(ݗ�d��a
?I��1�Z��Z����i��_P7GZ˫������f�d��b�e?_�7Lf}�ω��e�cygs�He�����0�[=��%t*���[ͶW�U`�)�A�bNl��f�	j**a�\�/��?5Fy�� `��� �Qd�{Nx"�j����*�(�w4�����eZZڞ�·�+�V�l���}/�H;�#�0q��Y�^*Y2�b�������$��)2��ͅ�����S�Ut�#�sHL�9���t�$�59�B�?3iл�.�ؙ~|mc糋�OcU������{���и���+H�t��|v�>s�����{��moKk��v�d��	������nS�.�HKt)��"��_�U)��ϥ��-TvR��,%/�ە���]�}�HUM��M��㥼���g���]Xs_܊�����6���T�Тd�(}�5&�뛳W�����E�8�Zm�ʑ}��Mo�te�2�+dnnn�[Ei�|:�Ne�c�����l�U�Ŏ��%�I��n-M���G��G���ɡ[��!��������?H�1��݊(�h
���LB�dm5)y'�93eI3%Azy���oJ��Klj��-��y'��``gVp�<�u�����h8�:򣣣��~Ł\�[�v��ǡ_է���Ȭ��h���ҟ:>KOK�-�}�@�����Pf9RU��5֭Z��D���fY�r\���%%���ݧ�]���t`Q�{�D+̓�`im�>�~���`)�.��v8����5�qf]���<<3��a���@��*8>��
g�*��
?Kn� ��������s��� ������l���n���fG�5�n��:/�vM^��Nmk [�f�;�aamͫ�|[ ���/�0�R700���Ǐ�^?��)��t��Id[�i�T&�r|�]^^�	����ӓ:Ĺf�_PxiY�7��C��0��>��=N����ս�U��HgMx���G�А.�v�4lgk4�^{�,0����4�G �4ܦ�M���N%�-�K�7�pss���h3�"�G|r��$%\k����-�4
MC7�|�^\T��6��<�b�(�w��G��<��#��e^�䊶��U��
a�'΢�II��=sj`�*�t ���q_���ɽ�uK�`�jwlצbm�~���c��M��+�k��)�Dsm����
��� ��A����	���)�H��E��`ɗp�Z�+��q����XetkS�|l��X jL*��ÖUTl����RvǣX���h��^�%����dB,�}��@Q[��-�[b�	,{b#o.�S�'�	��L�i-�
ff�HF�c���cY������I{36&f�W��|{}�uX7������FE��f�:"U��WH�Z]�G�g�#M!5vMz�3Q��E���5Eǌ��Ȅ�G�^�QG[� "O�j<�7��ͮ��G[�;�چ5�H���:M�� Ш��b{�5�`n��� ��*D:(I�ƶ��mt0�;eF���3���z���;�;~fffT�+�A��I�J���A[ZK�D^ˈ�oޠFA�N�t�X�����v��E�Ӽe�Q�h%0�c�qp-Z���C���*��D�(����z��c���;�t5��нV��~��l÷��n����P��yxD�Eo��}a����p*�@yx����&A]��e޻hБ��r�:á�r�ę���>'s��%��c�8��q�N��@�֣5z��$w񣎋��J,���͵{p0{w{�t�@���瑖*��PڀnW�\��'��c��4�:�%�4�ЉJA����� ��&w�F2R=��x���o���ϙ?0�y-��,�""� l9���xyyiZ|�JM�_�3��ǣ~������v���8��uj���U�a�D*�ET�M���|��&0H�mZ�����&��n��+���d矙�P"$/n����SQR
vww?u�hwWWrPP�����~���h1�@���䦧�wōQ�Z|��AG�ׯ_h녅��!��Ϣ�k�J����d���żݫ
��:���7t�-}=�/�(2G}����tѭZky��W�b�X.��:�%��y�����yP���zi-X���iޕf��?��k�����/�-�u��m�=)HI��߄mmm�X�}˄�f�Jݪ�A`�ٕo�z�GJ�l�����J���P�mKCG0��]뚼����R�!�,(sm�<B!rr���&oO����"#1���9�f˓/c4��N�L�zmgN�=�C��Syn�0�S[m:sM7#=�{���>~t����p{kk�L�C�@t�$vif����5�P�{`�B����0v��������U��D�S�%1�R�fff-���u�Dc�U�v///4ѳ���]��6ף��6�|����r��4jv�$���>�^��D�hvnnAAAY%�ڵQ��ō�����/S��na1�'�ihD�b&��^��]3 m�!���IHHx~9���W�UG��%��015m�7\�-Y��>x�`�7��(2RR�y�a�Gh1ry��9w�˟]oT�Ș�]ܸ��:�+��4�qH|�W�?�B/[*<sb��)�ᒧ<����۽Ҷ�pH�^mb;J�2P��N`����WZZZ�qUOx�! [u�S��$Yݦ8}ɦ�Q�������� -Y��}yo�x�ӿ��7�ʊH����bq�����#f�N
���
j
����U������>J)���☃��c�P,����*D��^y���F^�5�I��ˮ�'�P���c���)���3E�����v�����K���cގ�D�fx������2���4��9���v��!�5
�8����1z�|�X�Ec��& ��%�����-�X����S]BTC��I�:����%��Ss�����5�v����t%WP�^��a��҉��1z_��jɴ}��������@*775�s`jjF�����'�sCF�n��\�e���!�x���A��]~�!��,�R���="
z'���η;̤��u �			����NCOb���]?U�%��44H��	��Ul>ԉJ���������(�-.,gR��GO&������G`��>�������G���:;�����C���]]zM��\�9�B� i�S� ? j���Q;��_��knn�m���P�щ�w����7��r}���TrJ)%[�҂l���c+�$d��cg0T��+�e;Q��a�CB�e,��e�ih���~�������ߟ_��9�����گ�u���<x���j X�d��G^���v����A����X����}M@gcv~��(�����碬#k����je&&&��>�e y��dY���,��4}#�>�
[�������I��&1c4�p�[�'
U���`|W�i���^Q'�2~4����_eL�=V��z0�\�7�*�XRW��є�N5�H5M���V̊Tބ
?tŢd��;��|���8���a'�3K��{�G4%7��B̺@D二��T��"��+�y�"h  �ShQt�7�ʉ�X[q�_**d�w��A1�0�_@�g췻F���� �Cߪɳ����8���ѝ�@�?�n��~�z�ȭN(P{�}���<�;��/����$��ʰ����1�I��V���f��m��Ƴ�|�N����������9�A|�Y��K��O���Q��.��m��Ł4B~"���������������N�=h��7�;�/��3�����O�HA��� ��#�]�شri��P�5�i�*�� �#j�Mڪ�3�=WN�}S�J�2u
��q�$	���̌K��͗��+��V���+���\�` ���r�;�Q�������"B
dD�4v�KA}�P	@�ni������������i�j8�P>־gb�ϙ��Wb��� �����~���������N�e[~"�(��Z��тY3�q�ؾ&|%�����~/hOk���1�ù���8}�ׯ@�<%ǅ���x����*t��~�F �d��7?��u{�����0X���v�f�H�n��'��>�:`F�� �`:����,���4}.e5�ٞ�{~Z>�����C{��������`���8W���� 91ӪL���b�x~�^FY����%$:���,����|#�J^�D��fR&۟�<���u��Ι?0:�ݖ_������tF|sT�kh��\��A^��=󈲽��?��fdB]�t;���M�<�P#դ��&���i֠���>R���q���1����i
d�MR�"�T3��HLO�<��v�w�0�Ӏ���>�=xT�s�088H�~	��D&�}4rO�����2Ȟ�>����o�F&I������pAHl�^R��o�u�Z�\�'�ގ�) ?C�Zn� MPo�@�m�����cS�s�\P��y���-���P2��j��ݲ�N�O����k鰝��v��emCR�"��P`��b/}��0>������@qv1w[��9F�O���~o�����%	?
�O���A��uws����Z��|��@�4	�3/!�I�·��T�N����;Q�&��nF:��sKK���]r������ �x�s[[LӘ60�#?r'� ��LMA�B����{ol�m���4�a�{�=9������$t�����~�h����_FrX?�C���S������>��G����u�%¼~Ѣ;��vw���y%���8>�=�N-9�SZT°���C�7�R��Ȯ�|��h��j\}��z���>����͘�׸�
;/<���H�I�-�(|&3�f�-��V��-�Vv߳ո��	V�̘z'��=���y�`�·�����#���H�駩R+��`,�Q�{�A��%�3Ie�X�y����MS���+F�x<�}�����ƁkWM�4��\n"�k��Z�h��QׯQ�`bS��+	F*�+p�x��Z�?���?Z�A���H��M�Q�J�X�*�b/
��nb�[W����zE�0�V=�F���������ARCV,v�oD1��Y�H�#a��G1]��
YK^Ji�j#������_�1?�U��%�U��O)��z=�I�I[.`�}a�#`^�ךaJǽ��Mn��ϩ��uO
�*0�[�����z`s����E5�:����Р:~���uO��_})��L���ǒ�݆h(�^-��f�	��Z������gw�Ag�����k?�޲ί�X��7÷~ċ�_&�,V���"ی���{?YH,尒z���S1|s&A3��������ei*���) �.s��h;N�"x���ӭ^�N�P[���7��o���KZT YL����:���(�V�BT���WE��z�(�Γ_���y�o�~�XT�E�UY//�AG)�W�a�io�h���dU���B��7+�t�Gu�ե��H�e�3�͵u \+��?��`�֏}����u��=�au5�l	^!���3��a\ډ�������ha��oo5n4�@�
g�� �N6GV�r���K�}"�3sV�f�A\�g�a�Q��H�=dܽ���P0Q츁"�f��V�=n�a�Lz�@�n�'�C�(L��=+��"Dv�x���vSS�+�Td�ujbÝj���/�'���+dg�����?[��AG���˥w�JgC5������IJ��\�j� �+	.I�w�>qS?ǜx�ӒSQ���-	��.n
݄'#�X��({W�N��몳�E4��î<��:)�3P�H��%�-6�[x���[�"����������H�
��2�����2F�5����KO�)^���1�\�a�縢�9�O$/�����O�s�ݸ�M(9��F��:��z�=�x�C~-e��S�6��y�_�舡=e�D��%�964����٦��9I�0���.�����J>�4-��a:��Dd��dB���<ϴ�+V�,<A�I��I�$��\5���M�=� >3P��;@�,�ǎ�t�8(��[��bS,�r�s�|���o�k��6Bk�	��_����_�~���7���5��P�j��/��k"Z���ò����
��g����;�ad��MY3r?bF��m����lb�St�	���AA�J��2jK�qϒ�ױi�I��G����	���vu����4�ڝӗ�c��4Χ:�[+�T�Y������7"}�O6/�s:�ɥ�Z0x�Q5��ۯ�'<K:�"}�'%o�8��d�#�G}"�7ʚ�`���{Wk�~�:*��8е[�_��2Ο����(�$)kڬ*]��2�Mc�r"4XP뭭�윪?��W��&�ýd�^������^[��$M�C�$����y��QOa4Y�L�{9���~�>����u'�";[�)���r@�{?0��]�>X^&�m���W�y���O����-��m�~��*JG��M��'��1���%^��α���u�:_�(�^uA҅Ԁ�u��ن�E^��7Tv���(��pCJ8�9���r�%g�����D���1[D6�Ce��+���OOg�"ʆ�p7�r�?u`��2��a�	�ϊ;:���g������f9~Ӧnc�_�cY%	s��V�r�rڥ!�Ǌ�jjj���Ńg����@o뭞�g"\� ��"-k;����춈T���a����N�ju<W��݃t�xp����ͳW� iCD�Y=dTc�q��Ey���tm��nkqH�O�ؿ���:{ pUF'=���T���Tn��9%��[�LZm��,�	�!���՘��/����
Q�R���8�&AR��X�ܱ��Jq�����Հ	H1G���M�\XU�O҃�I5��F+�`o@Lx�@��?hh��Y\n�nNA���V�k�	�-kz�����O��w?!���?Q4=q=�$S-��v��`Aw�٨�� �6{ޡ{p�TS��m`an`�~4���R��]���*�2���Wd���T����զ�:������m�3}?���_/� ص�{G���=1�������VR���l�4�D�M��y+�VS>���5M�|��jV�����b�O��=< �e�kC�qE���V�B4e}=�����z�7��υ65N�i�WB̈́s-Eӿ�t��"+NxP�DP��o�o�;�i��ۊ�Z�n��*`�Lwb $�%�:�/� ��d�Ng��j'��,��m#�e�A9�͸g�5�{�VU�����J�yEx�7:��1� ��r���9')L���*&��@� ���po��н�E�{�Z5�Fv%fV�����Г�������M�����c[�OQ��v�`<H�����8E�k䣫�c�y�6�(> ,�
L�NAE��[���Q�y_����O��6���PWg�\�yc���9�H��O4=��V��R����W-��R
��4(���G@�/|� �7B8�@A���%Z
.�)�3��&�)�4�Z$�����z��e��isj� ]�<�{�p�P�>�aMco�����#*�riV��ke���q	��&� t���^�VHI�N9J�81�"<�K��K/-�lo�V �R|��9�<���M?uEYm[����DH��>������}���:CQ��+׬��3�& >
��)�{�:��S�@�r{�F��aZ���2��+4����}���	g�t�1��ʧ2���^Zs�tgOsP�>o�N(F˘�v��ZO���H�'p����YT�V����C���.hm���s�N�.a[���3�mG�qA����\# zh�D�Bs�Xg�1�:x���'�]6'��ؾ�O�C0�:b-?{Ƌ�vvx��*�S��O���Ԩ�.�ʺ��_�F��0�l�%f��R�n�XX�v�o ��q��Gkǿ/zߎv�H�%e";�	�\5+6��!k(p�j�^�j��KF&X=Z��h����L1ͻ����\��@���h$¦S�I\���Xҷ�1��?c�Bg��&���j��w�@�Ϋ��a�͞�3:\k��󍢅m��X��6{OB��`��Kl���`���k�W�r���5Ju���B�z�	�?iV�"��"�i�T�7U{q���~��ۦ���h��A2��g�u�v��)�w,�l��9�Ϻ���7y^)�������ƺE��;�;$_�=���<-�`�.o`��k|�:?��s��"�h�A���j �|j�Vr�Џ����;p[&Ŧ8��*X��c{郰T�fb8�5@�;�+N-M��7e���Ռ^����ǲ��T�#�����<�4��|�Ta�n��Ŝ�s|��l.��Ԑs!>_si��36��qY�_�6>7�ѱ�d��Xl�͈���;6L�
7�_�AD|d��ʱ��%_�1b��e��Վ�{�cD�,�'ŪQ�|�g���.�{�ZI���d�eIj��A��E�����35�4�+����a��[[HZ[�g�A2�> ���o<�*;;�w4b�C�5�xd�f����,���s�ֻ	���6`��m'O�e"̒e��$0���5��SV �o������hn�j(��Zfٌ�(M��.�~h�D�ѳw߷ P�I���Ċ���}''�@M�t��� 0FF��oU�uu,l� U`�WHC*]�IT���MH5�{/�u�BM�g��8���_�|�����;(&��Nn����-��M�ĳ�]���@qpy��D���.�[]���׎QxKUߕ���s��E�T��t���p�@�3@ze�v��X�O�˛�j�ۺ�[����=���}���;�_�&Zvc�Wx��}�\�[�@==�c��TR:�jf�rZty��³�X�r��p46(I v10�b��K���1abi�����3����Aj�Մ,/�b��XޱRW�+��e2�K\|���e�_�u������d�*�$ގ�P��ď�-�,,��i �/��-4�"L��V��+'�U��B�oxS�w����S���u������0���O_Z�%̓��8T�9[�􃺢�0�S5?�/9���T�M�V� �q�B��햙�:�������5*4�}Nmh�2�=��̐K�q�-��9�&����{���m��@��'ĵ��EmQ�c���k�s�-Mzl��y����,H�VP.���r�E���� C.0ҰC��0rE�w6�����s�x�nY-����}����
���e2��@����~zu
����|S_QS�Ɯ�}v� �����ȁ�K-eYn�ؚ ���a�M/��Ըi�w����R  �'��K�=)&'����_��Á��A����V��&g/�^7�$}ȍ�j���;ѭa�{�)�S1QQN?����^���� e�$����||j�a-�1��K�v�i7E�k\'<:�#�p!vI�}�ؙa[N����:��
��8P�;�,�b.�QIi�Œ~2�5Zu���lq+V��3��:�#O=yg=�<W���Fsz16+n�n �3���6SR�iw����`\�	�6a41��Jfffy^#W*7��[t9�|H�UH�~����9vc�<�/U!Ä��C��N������A{/ڄ��/��D+|�gdG�ٗ����5e㪮��b��	,�j<m;���b���_�(�\%���du1hŗ $�?�:�GC��Ś���k��f���:)s�*WxU�9!�h|�~�7�Z��>��sm��PQ�S�W�]�a�d0����K:���I���c�vL�JA�ۮà{]sGĢzi:ۯ���;��� 8T�W�:����4����ˏY��.�g�K��U��r�ZA� xI(J`��%�˿�/�����qd�
��5�k�"}�_n�6*<��>�`S����	��]N�:+Nц��j�����U�(����*3��h�����QHF�p�c����]�E�0@�D�6��v��P
UnD2�ǁQ����{�l�03��-kZ}!l�wޣ
�3��0S��2���/株��01��v�������4�`ii���N��v��sv�}���
���
������bP1�)�3!ԗ_Ѓ�U�@Y�ʛ�D�S���ن���?��S�����y%'����� �ؗ�8ox�NtnJ&l�AF�0~��*�r�b���� id�ݍ������l	U�D��) ��F�Ot����&HsaEG`����,ֺ�,L�/�� �Ǫ&|���\�=FW7�x ��o��} Z�{	Dz����SF�H�����/���Մ!G;��ϟmW�ʆ{�+{�Q�	 �o+��Jy+F_�׮�c���J�mەd�ۍ�
������O�N�������G>�ؐ���7�j`���&j �! KPW���Y|d���٨x�����$a;`<|�/�e-�� ���ы��>.R��~L���/^��j*p��	t�!�6�َ�Z���] ���C\�R���ҎG>�?�@�1	�TYu���jX���d(tf���"�K(�ّ�Ӵ.�>�8+��"X�N�&F��V��7�����FqWɢ����ߝ��:��~Z�8�KZ�����uʬuKȜ@#y����,ވ����lթ�6WT!�嗮#��G)�}�q`/'�`���b�YE��xGU�B���H��3��[A����I��,�_gB����it�m�U�z?�� đV�\4����|l@6_	Od"�_Z��b��5����s��'W�=ի2P���]�3�/r��j������׋�h��Osv`�zXw�ؖ7r.� T�������BL�.m����hv�h���ߍ���HJ���I��,Sӗ!��eQ�D��wDض-5��n��Q��Y�\�{���Ec[�ÏL���n���f!�/��Q�	F�[/�����0=2���`]�3��_��c�bP�a�E��u3��V��"�:��$_���|�����S%x�j:ō�g�h��nmK�l{Ǣ�������GrL��'J 	�C�(���Y<N}�af����+�b�c�C�J�G����m痍��n���=Hd�ho�D���	J�ve���S�х��ڤN�*�MAl�Nu��h��=�$ �u���*�Yf���y&IKt�VZ���Z��KDHћ���R���ă�y��Io� �}��zI���7o��1�'V���Su�I<�Ӏ,�LwN��z����o+�^��j�o<�y��d�+֮Z�c6؎���Q�}ؕ	����9�9%!H��W*o�F��=[Vb�`ނ�b.��tU�����9��vN�Z�c���^$�o45֢�>w�b�K�����\��j�\&�m���PSJ|��>��8f���74l���҃�!��Z��«5c�|���������2�lYd�ε���ot\F�8�����3f+���kM�f�������N�6UD?��#|��d�:,�xz� r�ݦo��ʬ$�-?1^I�����E	),��8�X,��5��I����a����"��3?!�V���0k��ノ��������z���)�o[W1���.^��m����H'�bF$ot*n���L�K�$��x�ȭ�(�x�Q�����B,�"T����w�:"P�PK���J�R�הZ[�@1�ܼ� &~��Nm�o��R��[�3�(����TĦ��Ph��C���۪|��E�	a�f� m.��� ρ|c.�v�9K�S<0�XH1���B����\�%N�����ޭ�ݰ�c~��Ʌ�Y�-d���U�,)bk9�F͇�nES�D���L_`��MYV��������Y���r�n"�s�v��Q{��7W��T���ێ2�-�I�Q؛t��.���#!t�-�B�3y�;��aQ�7g	�g�6݀�՚�����&-q1�����V�HKzZU��)̆~����GEб�Ww��~�ƹ�]
�	}x��-�ly}R��я�MGS@�7z�G5B��>ڂ�[*+�ŬO,�6)з���A������w���d��������Lom�x�W3���$_�P/�nyѾ�-�Wxu���ں�$(�d5z�o�S�▆������wz���Ǩc��v#����S�	H��� �[��&XR��"���\=�V���-��N����ݓBwr vU��0H�)޷�}�#���O�?2�W�^%vXK���'�u�s4�2����Ϟd:O/s)AO�{b�$Է���Ej`�Lh�����O����z$�HYZ~��B|�i��?7�sf�;렜����iN�]��u~j�u�A�]��f�s���z�Ӻ���T��aO__��?�h�ÎsF�ݤA��2Q���L���������r%�����S6���>S`��ȍ�c�&���G���1۰[��lگ7�����ˑP��aU�p���{��N�k���c�ڤ~��O�������<�69(0�����j�"W���Un�/��i7.���0��i�f�o���?h�)@RX�r��nf���o�W��� �^������d{Y�.#"\7��c�����[z7�g��C;c,��<��=�?d����"���}�8�!]�~�+6鹎tr_Q�M���y��]Xz��Z@S�
��Ǧ�Xz�?"�ǰ>-F� ����ײ��"�2�`ۥ�}��q�QJ�ǟ����(�ӄ���1l�׈H����%�����W�jcga�B�zn^^I�ݮ6ܩzO�<�y~�1Θ=���I�~�#��ǉ\i^�>�+H���Ҏ�'>�{v	�&mVw7l߲�+�yt��x�5�TB ���#s��VGF�n-�:�1���)7Y���{O�P��>,,�?v3PF~��y�v�q9;�
����H�����z��!q�'��ɷZ����kτ����pV܈BŠ�ϵ�tK�ڞ*⠚�%��!���?���6MG�n[��`$�b�`���&N��܍/��iu�\�cF����W�����&��a������z =��5�_Z���43�֏��䢎�=�HJf�D,���ׯ�k[�j�v�;%�r��-Y�jA@�,iZ���8�����>n e��9�z=�aN�����u��B���Ri=��d������f.f�ݏ��.9�&� 2�Ҥ���M�K���ESE��‍�x���rO롚� �t�ߜ���c�k_���wJ���@S��I�iii�mSjE�ǯhn<���!�R�W�1Y�ܧp�Wc?�z8%0H�]���-�'Fk���R�DV%��� [�'��<��}n���E��턗S��V�66�V�X�=�5�y^�_����4�?�jl���>5s<X����Z˳�u�Z鿔�~�}�R�#���;"ECX"���u5��겚E�s+.L=iL�
�u�\r0� �dW�גם���x�(�y���R�n�Q�wA�-����kJuI=�z M-�����k��MlD�nͫu�{����QDF�Mq��'L�WX��jIb�Q���fKDU�4���llɡ�퀹 H�s������Ǡ���ߠ$��B2�"x�>㳓UWV^o�2} ��@�������&��eU),��9ˀ���������.��YX��,[�b�W�ͱ ;���@�|����!c*Ȗ��0��c�k��x�Ё��x{�۩<\����S�����2XX���������ǭ�?����q�d�����3�o�0s��s��-�73>���S5�g��j�h��7��������B�7��W�Qc��nݬ ���y<d������� +�K��i�\�V�4��[d�U���Rk���/{fZ�]-��Ƅ�.嘤�zg4b�CR����U+~��Pb���Z�A ��,�`l��m����E��{���t0x���QF��I�T�.������� B��m�D ��58��;��i��"��]J���qt�ĐSԎA�]W0z�{y\|o<�c��\�pPt	j��6�]��������z�,�ǻJ����yKwww5^��\�<e��rn��l3�Q	3�����}�>��i����ܒ�AL�Ǐ��rsU��_Ѭ��^>�sSXq�z��1?R�Yh���[�0��I&N��A�v�Kn�M���rzz�����	�����js�Q��Z����a$�mm�C�8�x�"�3X��ٕ��� 
�P��q*�I6�QSSCq�X���~땤�>GHG�J������ �V�����^�
���ch\$5G���뒝
��y�g��[�}q�䋛�f�@�Í�@�h��X�4*�+��+,*:���q��@�j:f����1}4�/���[���|�U�*��X����~���0�[�؜%����j�t��KU.s{U�^�%I{��f�T��w{��7m����la�4��ö����w���+1�p����>d��:ImÌ��5�}�Yq�a��^�O����_�z�;��=�x���+R迵�iqċlc��������Ԍu���#jK7_T'}Z!'�.|��+�J!�7�$�r��䤥��$�%�-k���( 	���d���V�5%��f?⬄�:���G'�D/o�5�_8�x�r��4ܱ�����eK�^�v���y��33�:�T�?5��{,1/�ޓ�U	�Y�����Z;
��3�����E���-!%%®���Pm��Vg��B������I�½���s��q��^Ï^���H.���P����o��g�Gp�q		!����ʳ��E���� �⎉IXII�3J�4�ђ.v�k��қ��d��(�rK�_2ه��o��*Q�Sl�0x�����i���$�R�DZ�U�V���RE�{�+��V�Z��v>���l������ܭ5�`�3B�q,�z�w �,�Ҋ}�7��L���OB������75�pD]-�y����?��a-�MB����\�g�m�4�gI���n4�*����=���ZZZ.(*�uvvfe�ɷ��ի�Y0�J�s�����u�oM9eT���f���-�����a�{$y�Y��L�:�1�o�%�Ւ�Xl˦��[��Z�́y���/G#?Ǵ���ې>�k����#�$�g20������Y��O]���a�
'�2�w�^x(��S+�������Q+Q���,�|Z�d������8pk�L�s뻓&4Nf+�9�}A���E��*�8��"j���ot3c�8��r���%U���e��Q�U�Q�JSMr��8�{��e킄�QoB+mϞC|v���32�Ԑ��O�d�����2�6L4Ѽ�ƻ�ok�~֑�#��'���߰��7��WHZ�c\+�4��|,ޤ�,� &eڇ���ҚӶ-1ȱ,����|�ԭn�y�dV���7��1+JAOO���]����<OʊJ��Ɩ��Չ�y���z6#�����sc��n�q�7u�ͦ���+É�p�+x恻~~�D����A� !�+�: �w��w���&.��M��,�<{� N ��˗/�զZpZ-��oa�˷�S��skAc8���U8#��~1
���.q��%'�C�K�og_;4,|kq29��=����rs�M��3�R�<?/�fh�s��l�c[ˣ:$
����@���>��"bb� s�r��Wa���/�)����!CE2w�0HU�@^haOv���Q�����-�Av�¬&-+n�K8;:_�����NEܻwO�={6��N%y2˖��i�C~a�s,ek�v�.W��
�Y��ab����W�6��3�r���T磤6b�C$�}�&a�G�x�}���!�ys���h+�$��Q��bά���j~�Q���f^H-��. I޽{�q}���a�K\ ��j����w��o:�M)����C�a����_��	�T#�b�%䖏�}1�=Ck"�=/���������bG����3Jv[^�3�zb'��o߾��G;*D��85��#��&'�4����0�g�<�u�v�����+,,R��4Ѿ��vN�F�pt���`��O bW�����Qa`@����rc�4�8ʅ����
 ���Ĩh��ZP@��NV�f�m,���퉩�ߪź���G���^#��/�ﺪ�g�t �ou	�� �\���E�:��f�x21�7Pbh9��7������+[H��z��n���gj���u��n�������W�C��FoAQ0�aÐ�k�SnhÐ���la�QHH�}�8c��P����ʞ����N���8�AMQ��S��z�W-��x}��.���ﴚ8��}������������Z$A��xǻ���a�d�Բ-�/�R�e~�>��X�5�]���A2S7X�������E,>�aq�-+LB<�=����侒҆��������6��F�9��) Yl�N��d>X�هr����:/<�BO�Z᪜���/Y�E�D���� �jQ� �x�&v�B��ꞞPc��I�:���}�T+ܭ�L��3����<p0)���55Νw8�� �+ck���j**�@t� R������,GH� �}� � T8_���]轠����"�����%C4�da�{0z�m�q,���aPJS5�e���v%�gW�ΦzaU7���A%���3۱��&#�/�J]T�P`Ϫ���X@����I�3�?h�J���3�d��ƈ�rť=��i�Xa�`j�2Ȧ ��`P�T>���'c��KROT���!����)~�$nhh����QF�<=���5���'�{������RG���qVV֔�,Tg߽����܇'L�����>eq�߆?��%70�w\�e�~)έ>9���N����R����iQ^6I����qhC��k����(��F��z��Y:9fۚ����l�݂F��q����<LLL��ߟvc�ݵ˳Q���N2l��[a�߳&i�?�OOO�+�p|NNN��o���"�CG���'����j��
L�6�m��EDE�+S�"-�@T#k�
�9��WD��&���5���߹� (̐��U^���8d Y�	�sf�>e���P��6+��TOl����`�.OUS�����?�Rj5q�@ � ��i~,����a��7��1��<iI�:�z�)��⒒n!�hT�·}�u��_�ߚZ�s`8�����E"@ �K�o�Be��گG����YQ��2�0y�jZ�Y2���G �D��d��T��k���֗5<�$h�#�{+k�qP�X�E<�Zl���a�XWGV��i��	o^����������v|��{=�H[uY豧A]:��w�ʦ�j�Y*��O�t�{�?�����9╈8�H�|D���=X�7/��� ��֯�� ��[��� �_C���w����A���B�u�ss_����n������Dm��]�[�ћ�4ջ�z�I��^�4�V�i��?�����u�cW�Ɩj��8;;�o� !Y8v�iz�ˀJmF�����ix��)��ut�uA]�\k�0_�&k���n5z|7�#�ڇb���w�xc_��%�\�R�o(.^�|�q]�5�$�6�;Ge}����y\T�n.{~:�Ԗ?_:��[<rDZ,���Ae	?0x�%�(�zV3E�GCC#�=<�ǁ�����# *1��f���6�\��tFJ�J�TMaZDs0ϗ��!þS�qI�Ͻ-��]g���-�f�f�h���>�?����|�j���Q����U�z�ɓ']��~�t5#��� �,�<��(�}1�O����;���<��7��Ж�OD�ߥ}8N���Ji���xd#GKj�������_���o��$�Z������'즁 �vu��J\N�8T9�����G^"Tk�[�kc����uR(�C9���eCG=&�g8-��%S��g�\_�ʂV���X&�4�>"�X�٘ά�?mm�|�)R�s�u8�X�^)]�Z����:�wC?眪��|���sȩT�SҞ��=?�Z\���<������Mc4�d2juZ�����S�����NP͜�q�RB��g�8�g-u�1#�^����\�Cc~���'2�(�[bh�����P#R�$�i���P��^�[�tV7�j82���I� �˪R�6HƋAeFf����?�mIþxB�R��IUO`� ������^�Ǉ��N�҂ZG���E���{����;�f�������^�H�G�'�������tɆY�ʛ.6ǂ�M�{k������+..v^�9ruVFӸ7/�r-�(t�W{2�imҸ#��q>�΃Y��U���ￇ��ݦ���dmi>��Q�]�h�@��l)�����5ӄ?���v�EMǎ�9�Z�͹��<� �Z����i���i�ֳi����'���ܠ�Qs%�à���=f��qy�|�$Pf��O,sYJ�����|v�O�����y��S���o�/e��OqWk�y8�0�mc���.�zs&���*�-
}H�p� -�ѣ�O����v5��W�J�{�=҃�q�y���pImw1� ���x3z2�'U�S�:Y�����/�kci|����Ȭhe��E��J�4m2+������v��tܶ�����R�Ԅ[�H#*�˼�q9lx9,.>��PwZ��U�_�&�r|�[�-�ٽ�0C;�n���иAGW��@��l��,D����]�'A�0c�㠼o��l6�[V��2�K�	v%\�x���Γ_����7�u�kY)�Y��69����#��1�ԧd�"B��"R�C�Mm���(5��b����*	���e$_|yV@@G���A���M�ɿ�k���}�4����~˖T�	]+� ���F��p*e�V�	Y.�R6�R��cKT��b,�Ĺ d	5�M��ZB��C���o����dC}+i -%k���l��j1�j�Xn=@�윗mH	uB-&@�aP���P
'LT�/���x���C���:@}pG�B~�P�L��d��6ķ.����j����u0aF��L�:7:\��7p�n.�D@��Č���զ���,g�M�w{4ÁW� uP;���e�xc�s��,��kk c�
�D).�R<"!!a�L����
��>#$f���/C��\��@u7�_Wv%��]�{�Z9>���C��t���tu�U$U,��t)c��~�>ǒ6Lt�����$���<k:Z,��YfNR�S�xz�1�u���I��9��M���(~"��t8\��}]��H7�u���9�^�A������r}�Qk���V�j��ҵk�5r��lWb�d������Ě��q@|��Y�����>\�f��'�(]��C�uکsp�
��dd��{�����*�G��D��������Llu�G�ŧ�R�_/n�(6о�Z�y��XXǴۭv����jP���ɞ{�F�+k+��{�Ng��6~R��@?��y�9�幊���ힸ�x���?_���Ԡ���
�L}���zs�z3��#a@���A��VIN֍/ʦ�s�T��-s2	�K�飣���4�S���w�� �`�����P)���&��;�1� 8@{��b��HD0Q�I���&6�E(T���{�Q�r	5�"3�o��������@;��t�����O�BV�ʹz��'���gW�7�T�r�,�$=��fiZ*��\��&M,�<�s��L_ĩ��V���r̷����O"wS$l�:��r����$�K,t�?�s��U)�Ǧ�Z�|zu4�v(0�@����Y���;�eW�4����9B�<������zM_Z,���ϧ���jJ�x]`$S�ql���1����-9(�%�LVg�����}?�23%o���Z����1����I��C��NS��=��-�
��s�y&���Jg��5�PNw0(h�t"?/ʃ@R$����5��Pf��!ⳃ{�X:Y.��� �ۥ��#|J$����O��X~�M�����:��qZG/�����6�.��d�������i2���nK�+;})����9�=�WF�m���hW�*n�$�w7��X�KY��֔K�K�nŮz��|�.u������l�ண��`�B����$��R;ڶA�� z��|[i���&�Q�{���&�)_X�# kF�a.�jI���XW��j{]ɝg�C8Vb7YdF�,�1����@P�F� ��vhVp�8\��-�k���#aW��8(�����q�n�X�IQ��A��V�H�Eq������ZN��'r_i�~؉c 7�6K���T�*i��p{{��l�0+}G����Vּݟ��� ���~cf��,J��ł�`�	�9�Q<L/�ޣ�(�	�ϟuwQ��$h@�=���l�V��s��z�P��r��|��������� -���
H'j^����j��>����k�8 �ɩ��/
w�K�%D��~u����0K-���F�{���gfz�������V���zO�;N�y�ː��n���(SS>�F�E?�[�H�����w���4�aM�y4ǁ�g�s��C�$����,mcvBLE^c <�JΣ��|k�i]6��a���д����u��2������{!�uq��>¿��!7�
��e�d��V� C/����$�"��7�g5�@�ǣLC����&t�zz-��}B�	������q6��a�|�E�E�_(w�5O��5}`�7.\�8�����$.Q��������OǪm��H����b���9�$s���ˆ���J��}���u����&G�E���޹}�������|���X X~}qx�e�Pf{��w9�
N7�!E��&��Z2�0��2i��j�}�"-��t�Z)��IF�������p�8��͉��8�U�9��<�1H�w����7�@iY9�k�Y`:�;ooR|}�C"p��������{��_�p�ۇ�:�9L�R{�)�'Ĳ)��sM���#Lf�Ч������0�M:��:�3c�����SV��ؼQ~�#?*CB(U�p�qߓ
�Z`�Q6Q�?�G�.�|�b�}h�ҜҼ(?�6D��W���`�r����b4t$e�+c�o߷5F�@�^��Xz?�>_�Yo�pgh&��4�'&���7��V*�QD
JY=T��{�5�� {�:?<�qV���l`���(>@$�Q)�V_�|�������X�T���elvP���/t����:UJ��pEɹ��u��������d2��{L*����Y�#"P?�.��I�C��_{YN�����[����9�&����㧠}U���o � ����POw�*n��0��4#˭��GmN�+�ph�h�aL���Ŷ�U[ĈJb@�X���a�C�?@�u����M�3�nt=�#�����#U��(��P�Ba���[N��Ү	��ܾ������R�S��n�4�M��k�Kǫ�o8KU�̲5�"�C]*@�$�g Ԫ��4=�'�"�^w�<�R��gT�C�=Xr^�񰁲G����@����t �钐��\#F�R����Hx�����XT.�������<̬�1�^�/Ԡ�!������5!}����T�>�@�����;*����G��/�%���PC�l��-~C6�ӂ���n6�4���h&��,c��{�U��>d����),-��0T�����nV����:����8` ���J+!ҍ�t(J����7b R���"�ҝ��|4�9G�}�13:�{��g����}	Wv�J�Ϲ���+G�r����Ε�z����9�[L,�:�]z7ތ���x`�(MZ�h9���(8�!�e�(Uړ�}����W��Y�̜ӷ�5�cF�CG��_�Ǧ�al��~���<_�ƌ��m�
���L�kf�z�<
%U��5����33d)|����"��2�e֓.��鋺�|4H.�7�t!Ρ}�I~�TSڇi����˼3s  ײ��*}E)wo���<��&L�	���+sg�=�����E���.G��.����@�C����>|����L���AQ�ڿ���ڽ�t������t����1
��0@2����i|.��T(�LޅM��p�'��*T���Xl�8_-z����:D�Ft�\�z!�yG3��q�c��˚���鎌6'���Ά��4G��^[=].�bJEW���ܟ�3�d�`����:Z��u���^@7��a��h�V
���s���̫I4O��B�++k�zEĉA����q�g%O�R��q-7��_J��S�o�#�P.~�"�t�i������F�ӛ�&����s�[�pI�>r���g0�x�
1�y"��%F�K���{������VY������2B�\���~Y(�X���>����W�����3��3(HI�+*�iJ�[bF�y�����J�=�n. c���<�����`��ݜ(�j&��YP�9�Uq�=�yDC�/cu�����-�g����]O4��'�_��q���@�a��?���xj�9qJP�i��$������E2x�#����?�B��H�n��@��i�&��8�'�?)c�b����{���q-�P�FѪr�����g7�QJH�}��D!�d���Ν`�`I�5�G��S���(-՛�<�U�����o�[�ń?���w�v��U��+�8�9%�}�{�Θ�/���|5���'t����s���[�C�Vo���#==��=��E��/'�_���@{����Ϲ�O��%EP�44
���S�^�P����X\!�"���}�S��?Z�o�X�/��j���	�qs*֐���U��
`�?�f(c
�ӧC��8{X����p��L�	ǿݟح�?4]7l��$?��%�8=�&9�Ԙ������Z�I�Ac7'�c����w���{�A7"����Dߠ���� �*1�$�# �{�6�O�
)A�s�ǘ��F�!��o��Kmd�{���g�p$F���^��"�����T��+��Uǈ�X�O.w<��o�Fy��,�W�(B׍���mll��A]|'<m��w��P���Ǐ
�I~�eW�R��ZXK���w���$��|���ǯ�X<0r�����h�ې�#�F4G���ʥ1����k �#1��q;?W�I��?mF��H�����vPZV������叼���K�����8$.�LMM�_��^�3'~]�.X���㩮���K���iD������S�.��1 t�Ä����x�?�(�_�O4|r	��,/yb��`l 2�W�
�g&��E�g�_�H����_�;X1�b m�Տ��~b��0)ݥ�/���L�)�$�	����'�[NB�ĔB�����,[t)f���C2L@��4p1B�<x�_�����w3��S��vs���IT{�[ۻ9}���g>������s񧶫wmd󢪼������h|��A*�}
Q��XUtH*�K�Li����ܿN��K�v9�b�zW�"��^�g��{Ebl�,�Ѷ�[p�����h{���Ύ=�?�C6� �k�`��)�B�3��X�}��������7���w��%���c�|�����:�_�׎MQ긏��5��7g�h����*��}��>�^�3���H�h��-�S�d��"���X��LT����D! ��E#�dʛ?�T�[i�Y�rE؞��Nl���ݪ��^��|f��k�	gs�U#ມ���Q{Os*��mg�NJ�_!a�A䤥?M��= ��qΣ5�z�bh�?��>M-�U
������������\=�@m�(���mQ�����`dP%��~|"jƊ;��V���<+�yo_Q�l�����F���Q����.����s|���e�r�	o���n?������'8�
�=�q^ws�.)y�S��O���Y�p�1I�*X��@�������ޞ%V4~Ś6ڤ�rY|2�5PK{z�Zm,��!�w�����:�9e6�<�.'�ٳ���W�:=4K����Q1���%K[�AE���0A��z�,��)��+��j˥��hnUUU7n��˥)RN�aS=r�p#?r:�d�
������ně��ρ�LLL�8���������dq�[�U��x3ʈ��ܨ[��|��iT('p:��mjc�_i��{�V��U�:��pǶ�WL���򮯔Ebl	~�c�W��L����".O|����aC�3C��I�yR��;�_�ʲhr��k5�iB(4�6�������I��g~�����ʂ�1��S���7���ta��t�X�q)|ic��n�=���Fd��Բ
#��݋��*�)�L��7�^Bң���cD�w��L�"o j�*��bF���t��Ͼ{�̿ŕ=.pl�a�Xm�i0���XNt���{0���|~ �7�j�	T XB�g��4��a��(ț=^�<>rx�ݰeP�?�����.�����N�J��
�ɝ�X�J5@a�w1�b�ZI�O�{����}QJ��������'�$���f�N�B�Np���������9���-�c�Zr �l�y�ZG�E$����eZ�tdCD:W����-v�!k?t�jWFJ��葹��L�C��$�ɽ,#ls0-l<FH׀�N{W�@V���:�2]�{m���
9��]�v_l��NU__�(ie,�����20v�]>�K�O���o�?�g�`�,�waa��z߮AtX��>�{.[[Z�[Y�����w|���%�>8�F2Q!~K�6=V�˭�W,��Q������:���:�^T����NN����4�!�O2IXGI�u��k���]^�
Z}#���R�VG��R��d�f��Hd��"�o[��0��#/%��P��y�_�մ��h��}��h��w�R"��N�����e��S$l|��Ϟ4�k�bh���\��M��o3 �B�Ώ�(;�C��-Hi;[FY�ݴV��~����h�y�I4:�")!���B�&x�ɀ]d�(�Ӳȏ��k�9���h���Yɕ���^�K�Ofɳp�S�#�#��7v��;a$�T�q!q-��H�~Z�@	�W�U.o���,,��:�����=D���W������v���\���sєm X4ە�o�����ٹ鿊�� i �PY�����3�+/N'���t�j��J�	{���2��#" Q�~�����kR�Z��Ĝ���H"�H�U��]T�{�=����%���A�5��m��#��&��犯�� u��׀e#��~�I W��G�DA,�>�}2�����)?��%�3�om���npӚ�S��z�/�҂Q��P���.�󈈕o=O��FlĴ��)))����>�_�FI�(��)�&v�<�qɛ�[ct�wR�*M��_8>{�JM����|g��X�Y[a@i�W~���*I�r�k��el�>�Ks�+܊u�q,�d������"�V�ڤ^�'U6���#�D&~���৤�v�������DI��-VF���1�� tH�9��m6%��D�6�|��KA����+�,�İ���[R%���N�g=�>�O���T�PQ�3��!�)���b_�bRXU�v�r,��e+��^��h�PR�ET]YO*�!�w.r|��E1�#|�s��}�;���K1t"淬���R8o����9��d���ꧧ�א&�jpSiX�x"���n+�(�	ʫ��s���8�#����v&�t���#a�8:�x�%�<��<�R�1���ߌ��c�[���0��\��ؑ$�����R��� J��)�˲S|���A�ޤ}S)�)lon{x�e�\�=(C��S�9HĪX�A����w�L%ߤ��iܺ��l2�S�Zl�d��Y�1_8�Q�:�0�\���\	H ��f��� ��oVa�U��k����5`Mϙ����gi״��@^����1������q����p8U�^3V�7��|:;;o����3�By�~��{�����o޼a��!���M�6+9l}9�w�ŷ�H�"�Q���få-�tzS�e���:���0hw��D���	\?S��'Ί�'t5{[����6�nY^F�5p?��%2�&��T<;��z�D����RRo�H��?_���i�j��Jã����DF��xFr}�v{��~&T�0*�g/j�;���<\'A�V�e6�(|���S���6�����#i2,�F��Q<��ʿ�X�i88a���׀���
b�i������?����o߄.]�D5���<�|�aޚ�Z��=T���0��Mt��ė��_4�p����D�����&`�45���?�d���XU�	|OOO��(5�V�܏�������O(عקN�E�W9�V
(�4��ML�
���+����r|;m0<���O�Q��؛�;��Y"Q�pvHW/dB�`dI �Wq�S�V�94@�o�W��G�@��*`����oxXl����+,E�b`@b_�xTV	�N�1	��P��*���F��2�Zi�]���7�>�E����s�oܜ"��xԇ�f?����r���QP�6 Sz3�=cc�~�Ǣfb��?���5,,���4�4L�"������*Ww��;[�ݜ�V��,~�I���`(Jf�r12��/��x�v�Vo�M����^H�=U�P�Ѐ� �_��U���k�S+��G���$?���s���;m_xt4��.Uŏ���>>� p'7��� 8�e��	4Ng ���k�H����P�L�p$Vo?��l�������`��&Nߘ�	p����O0�b�1Kb����(I�`(�c�1������Z�Ͷ[�:���u�"2@v��,�%�������yˈ'_�%@�G�?�]�Q�!����\���E��F����i�Vg��@���"K���D+�n�xC+k�Jn�z0����y�]g��*�:@�;����֖>�I��~����4�Xy������a�(Z���[�ųE �uw�gT5�m��V�v� OO�yN�ֽ������mܝT4�˫S�Ẫ��5F$����pO�aD�X8�3�p.ΰP�z���e=Y�-�/�W/�h��0{?%9�,(����.�WE�Ҝ ���6	�K�v����Un��K���	�k�G�m�fp�a(�(V�0��2�M�g-��n#HͿ�3	��D��Ȼd`
@�8nL���]Z�"�����\'��+'tlw�a���� ���p�	����0�ӡeV��1cw�骒<�eJi���6����0���m�&�ݣ��k�R���t/��Ҫ	b�o@J�Wa֦����2.���b!��+S�����CN��ҳ�����>`�+�_�Q��7��'��PKM¶b���^ɿ65����$�U��b$P�vFن3�[aY#x�e���]��u^�d@��dɜ���rC�~�9���uK8�Ԣ�B��ۃ? >�7�.L]U�"��0Vy�dƓwKV�3�w^�m�%��%�NxCx9M�W-A���sJ�%c<�.��LG��Wp��WYۧ_	]=^-�>p�7oz� ��ng�cU�6��!~�&E�?��"��ɇ'�!w����Q=�0b6fĉ{&�y�������G��ἃ�>�آ׉)�T.�ۛ�ةÀ��ȝ�b���m����+/�2�*�`J��ư���҉10����^��T��#�溜�?�{4�;���4�|2��M4��x� �E���CL�2���� W֭)\w&0�� ν�8��O9��H��YXY��*!2������� �Mv������`��ݓ�h�ĉ
�k�Ô�Q�1�?���E��VI�,��������y���W8����2��k�M�l4,��Zx�e�w�C���es1NLG�����o�H�d'�b���
?]����S���.�;6�s ���i%*x"7̏dZZZ�O��DC�!u<L�,mÉ)����\\X�-$Ϫ<r�j?�F��ϣ�(2��DH\\��8�E3p����J��WC}9��CD�5"dg����O�������lBu���1��X�%�u�e�8�ʪ��y��vF���ʃ k����U��KFڌ)��K�ٴ���r�O�s'ФK���U����Q϶�p�g><<�p�Yu��<��O(��sh��	Ɏ/x�9�RѸ��krWýV��xyOV
nݓ�F�c��0�	Z���gFd H?�,5,�H1��چf�]�߉�ӽ�����FNL0(�YM��'�L�=F^T�;����ɨh��uN�K���h 3A!���e��)�4S�������)���/��%�$W�~av�u����xYu_����R�����vK	���'�Y�Ɵ�0��j�fU�F����tX�IJJR�;Y�R���V�IOS-G� H}��#�~}�0]57I������0ky��F~kkkA]-��
e�n�Q'��Y�y	���^�B{0M��� ����pvو}�᧱�D�T-̃�!�������f�_#�Oh�����(&Y��
�7p����z��������f��ҨG��!����
��ȡ<w΂M�Z�X�}Ç�Pz��HX�Dg��;���())Y�������T� @�@�-���)��� *����͘���)|��-ǧw�oPP �W��f�@H@�|����9��Zul>���I0��P�0iC	Gp8�k�Y@� !<cU��%U) ��s%����,,,��0�঩�j������<�W*�0h�GT���߹��Yu��m�T�,&ֲlS�~������մB�cxSvvۃ)s�#�����R�<S(��K?���Wa�--���ehs�Br,9�o�w�꾿���?�Y�y���XPR]�"���]QQ1e����w��q�>�������OᲚ'�wd�%�%��K�����_y���͹rIDk��0Ze��C�6��x�j��Hf�<�?p?�I䱻� ���/��u3�ݙ���^�J��!���iJ�۸i�25nJ�2� �G=i{�^�	!��zЄ�m�``?*�HR.�[Z��3�V��D���Nh;�	Ǚ�`˕⹺[��H�m�Io��l�9{6)�j��ȣ�<܂;>�F�yc�V��v�t���F��_�<K�#��Y��ȴ/]bs�ohL�gȀ���(�.[����35�f.��������!$	�PFn�{:�̻���isb�3���{�7��Z�"�S�N
�����V�py�_{uV��~g���Q��"!� S���8��~��s��e�M�ਊ���i��U�~��R�G;�h#<�x�ɽ�29�[>��-��� ��nh=���_R���!���	�!: y�~��0.�eve�B�u/Ӹ�9`f3̆v2��;p��O~�oyGu3�?�(�=.ג�D�� Ϋ*�~�������VF~k8k�y�ȝ굱�}�j���$��fpMܴq�dr/��9^ '0J�}FG��2�j�	���e
)5@d���-���\���]�?���u|����ˀ�T����LWɾ���byp�!\ R�]�.�[��{����d��O�za�`�)�=�2E�P^���x/&��5��gr�i��#�I��؆�������aY)))��K�d(�[L��if2M�(�G��z��R�z���<���$��[�l��%����Z/���l oT����8C��c�^�H�嫵��;���T�n���x�4�G�hJ�mzI+ĺJ�KU��J����+�*vΣi���ǔY���ˆ��ٗ�y���ck0�ҳ�IGf_�/%�,���hڔ}����?����D q��!���X2/"�6�:�˗.�<Sּ�%��8jhkk�-�.0#��s*+9cL�,AL����R��N jw �:���|��oŤ ��� у�%�}�� �niٿv��^��8�����5m��A�s���0p���Fq��;ڦk��o��@�M�=��T@�s}CR��A`�T��XyU����Ƚ��01U��7O��zS΋���u��?�Hk���\��D���� N��W/�ڢך+�ã�u�}w�+����>߮�%�3b��;ޔ�l|�`��=���R�`sӬr�����
�C�� �ϩ����x�4}+Wf�������gv�ni�0�&᎟Wm��'y��j��y٢��1�� H������#{ї	�y�VXJ9V�҆�5/
�G¡�W^�+E�p�N_a�u沟�}���`���))<����3#�c�)b�*����	hJ,Lz1�BY]4=�� ������1�����Bx��i{%
@�s��z���Ay%ͳ��耒!��4��[�+��[ևʶ���Rװ��;}JH��s������o,��
�<on_9O�iֲ)�+�ؔ���< .���I8�&�PY楫d��A��Yt'w�
�U�1���ܲ�˸����Z7�cH$�����$Akț�҈���P�O�K��4鳹ڽq�8.;'��?�/lߪ�g�<N׮�[��/iVBoV�@S(����Ė�������(�򞝶?���8�����!�-�?��=Z�MThdk�E���#���g��?�"��:hʪB��~~���_m�����K�5d^Y���Y��(c�B��<�ǵes$/Jܺ���HY��ٰ������<��w�+�`��fn̢�2ΊLSw�j9z�gEY�A���xO��k�,YL�F�9��� �Ɠ��.<�Zkۯ�0����l����ape���ͩk�\P�fCL����E"&ov�>=2]��	��������XmF�h가���)��T����ʅ�M��Z�����Y��*f�?�VW.)�/���&���W?��>��<��NO�潸r���5H.��|�m��2!�i�i%a���F��s'����l��u=��+��}��+x��0�x_�&ȟ#&66lf#����s�w�T쏬�u&��6�pq��װ��1D�����W^���m%���P��!Hax�RN����~�S��)�b��Uܸ�Q��0�f"��+7�@
�q�vC6A�ٿ��hּ���>K���Ę�yQ1� ��7vwJ���:��Ƿ���4v��)g�B�T�1*`t�/D�2�t���>a �[��E�h��sb������G��7϶FN!�h�PI�m�y��գ��:��.f��Y��������@��(��/9u{x 	y�s6�#�ݒ�h�{��g�����+x� ,� Atm ���i^��1����նaw|���L:}�W"94r�Jy��	����w·3�&?��vԾww���>Ё�N���h�>7UGb�_��o}Cp�S�F�s�g�:��~mr��x)6��&\vv�΍��=p�lӯ����>y���7xk��c�żnw��Mڦ>`~��/�:-\+���`v]��v�]�&V�ub��OM˄D��mU��n�aiI4=�æx؃ڒ^/}��o/ �_��h�A��	\Cǣ�h^�]n�����2!�7R����9;����H��4���T�.d_��� �R`�����l��8��B��m�z�]Cm�2�ڸ�0G�a�5���b ����k��.�Ԋ��YZd���	1�ǲ@ɺ���i�7���>C�",#��'q"78��_dn��aM	�F�G�>O�� �����HӰne����W�*4��o�GBr��l����������'� �HG��.>>��Ȫ+:(���P�.o-Z�q�%�t������Pa̝�I�;\���W�E�aְ�A6Y�!qDD�f��M2�yE��RXp�� o��$��fn_�*>������<4���e����h"Fz����������u�j�)��m� ��Cѽ���@{�M�(c��H��Ճ�հ�+�.P8��Č#⺤Dn%3O0:"�?2e�5G�9jO�9D`Zf��7�\iƩ@�ku�x-	)�.$��Nv��}�g������RˠQ����iF�ؐ�i��1^���
����������F������=�@����46�[8�E�����/�pp�����2{��*\9R�!w$n��>x]C �+%����-��OY�k"��b�X��"��ߚ
B11jB[]]W#���r��9�����A�
�:#�w�b3lv��Wc��dx7ZX�f39�_�br�Őz�G�v4��^�,��$1���0)�`�0�����x���>L�����5��� &��\�;�`P���~�D�ۓ�F<EEE'��l�Zdp4z�R�ee�7��Uz9�C�۴7��e3ca��0Hr5�u��ָl� P��m��G�0�%���	�־�ŭ���@��@`$��#��r��̤�$K�����*��Z���ȣ{Ye��Ɇ�3�n�jV0�$u���F`}sB�PR�D5���A]-c/W�7\e?�'�l�j��_��]��U��32��6~f�?��Ғ�A3(1!�)V�~�&t i��H.	���I/��c��؋��5]h=��;�D�a�����l�ƀ��B�s��>����i>R���lֳr�0���%���>��.)V�R�a`��J�6�����f����vK?�vU+�/|
�L�qʫ>ٝ^>�<ރ)8�sB~o_7K�%����#�^<�vq�#Iu҂��b��S�V+#�j,p�?�(< �͛�J�|y#�/��;��=r��oe'��Z���J�mkZ:��:��}�9jO	�ER;�_�N� �f��n�	;���w�>T��A_	�+6�mĴK��%�giJ����m�L�O�r��~va�1ypd������V���v<*	�p��<��f{7y+� j���cm�G��<[�M66��9vso�^�W���D?�`��N*�Y�{Y�C��0_�W_4�0�ܿUQQQU��<+c>V�e�󹴴�����#@M��-:�k��
�]�+78����_�0 VV�n�% AM
v|M̗�x�[Y�� E~��)��pOx`�iɩ�-��Уp!�q7�ug�e���jy6x?�d�b@�wc�Y��M&[��:iQ��se���&N������Cq<�܉q ��P�ȂY6zG��.V����!��?�˪��*�#"_��Y�H�,-X��������3���T�]x��P����L���] e�^�¯�Ў��YǭE�d�H���E�c�4�B����&6��`"]8���,����Ua��`�P�V΀9#��ŉR������I��a����Ax��t𦮮.�DN����U�v~tc��]g�9a,8 :9˞R
��)�9
^;�
t�j�5�NX 3��Q�&���1��d��Ru���'�����jb�@@&�%*�C���&h����}��_YC��1 �
��8������>֬���L�'Xsd��%و}0˶_�5A�_���B�}u���_�ឞ��ɂ>0�`�	���N�<T�<S�\I�S��3L�^t�^��d�E�CT��� p��,t��M'a�$�ŧS@U�4*,�#9��.���=��`+�J	j����˵O��T5����-�O=�����Wm�f��|��A�d��b a:�e{�G��2�Jp��

�#a�@R`�2]ϴ?�\��7��T2�P�:TȌ�S��ZԂ�#\��$g��i�S��'�e������2�NM�z�G�N�~�<��R^�tӠ�ׁ��B �}��+�1�<��do1�=�#�P���!�+��f��4�<ű�ű^�x$������/K;v`�����Z�@L�C�E�)�����	�%I����v'�$��k��⸀g��/�l1R�����+���*�zr���Hʻ���������!���� ���(z�}�Ԭ�@@@l��Z��a�g����rĶ�V�r�Wd_ê����'�0�44�'(0'�TO��h�����\��hS֖iV9�1(z���@.�j� �|�������*atΓ�����w%�1���������Ǉ@58߁_���<`m�a�&�J|щ�]��{�1"�|��(�m@�UX��w�ֳr���K�w��;�L R�(��B<Z	�e�q|a�%F�RE�'m�cb���W��jnG�ep���m�"���]�-�7s>�W����&%�>�{.Y�؂���keT�_�ɥ�=�pr�ʕ�$���6��g��Qѽ��SA�� �J'{��G��Η&'�x�^��R�Ղ�g^�ߺ��p[O(��W˴�$��U~!s~��)r$�v�n�������g�f��~�9w�F�������ѧ���e�`�-�[��c�Z�7\˝G�[�b�O���
��InOT���v�O`�����ٺ�#f��?QQ��P/�T�#t��q�\S�C�GL����?�ٮ�#�B"��'������5���4��~�ݻw�K��o9�!줦S��z�OU�V�fS����e�|_�2v�\�8.O7��m����@���~f�_����s��y*�_?&�w?3*�����$�Os Dn��(cl���Y��Ͱ��բ����m���x��+ ��6Px8/V/��%��^��%����A�[Ax��42��t0E1��>��3����v��f���ti��9��5o�{z`~�z$�䈬�����}?�VU�Ւ� ��}zZO���'�Z��}��r������e1��σfK.��N���	0��s��XI)�=+���ۛ���~w��R
��r_��
�!�$$��D���QPT|�ev���@�d�0��Er�'����b�w��4��������_��
���SZ�;����?��rr�z�o���J�c�2��P�RC���̱~�ve����K���Eq[��LOg��1�

�ҥ1kU�YvF+�$8����g�4��O�ӓ�Ѹ,�A7o�xR����}yE��mQ���$��О�;c����v�]|�ý��'��F�&�J�b�wcw���e16�"�������b�;n lc7_1Y�Yv��!�ub��ѩ��_����g�u}���/l��
I�b��b��j�Cz�=ꔚ����b�i�jbw.VLY9tI�l=������	�\����O|�^��"�z�*������^�(ѸM��Ǔ����ss��z��n���פe�=��k�����E4���e�M��r��<�;�Bq6��Hd�d0]5��Ƞ��7e�2����'�9�LG��͛7#�T2���n<3�\N׮��H��a0a�w�:D���tHk���<��岗��ewcn� a?�g|W�:eq�$(8�8g��*�K^^�CV�����g�epD:���S�u�x�`�]������N.��*�%��[�;�Z��Dw��K��Z�+�6���3G+!!����|�)��@H�������-nn�@�������9�����i�� ��p�O��d������~�;w��?I[('TE'+�i�z,����#�@�>>{{�Z��vϳ����C�� �@�����.#CVy9�y�a�W>�/9����Q��z	�ͬ��0Ad�\�Pi>X�]f��^�������9zwKMΧ@�!�Ԛ�4��}_��7��V�� 3����%�B�g�ࠠ�f��e��4�;kS��z��z��>4�[[����u�����!��ڊ��� s~y���jƪ�����À�G�}]GZ �X����&N����+Iҳ�����@ͫ�7>FG/#b�E�,z�J�H��񷓁�9\l-��HI=F�������&�S��|y�)���G�N�d-hKp2���G��`��������EN|�A!!��Dېރ�hQ*0�F�(�O�W�fS��,�Yٚ�m��E~d�JoL���k����+��.���|���	��B0r�=�q@��C����k��C�����?j�o���}�����=/-���{zp��F�zz{���ϰ��sYN��>��������Sw��Sa��l����*b6�M���?�� �/�_LS�RJ��&MݢXCa}����i_��yᐼ�B�^ɳgόLM��,��j;Qq����KI��`�#w��i	�]��TOh��~����06��Sw~��?x���D�����Cs��"��c)�i�;��bD�
���I���)_�0f���t�?����"����|��3�5.9����4cp�t$s15��Խ�L��O���m�� ��"���f�>�����%�P3�u�J�	Z�]�Q��09t���y�u{����АJ���E�}	���Z���=�ѹCȬ����X��-�Ѷh^ve;������ě�s������ױ�r�+�r��B�og�����������ք�\�����+���]�|Y\F��A `�Ց�)�X�߇��x�J+%�@~���/,��p�}-.++jo_��+�����ެ8���L߿'(�j^E<ztX� uV��ܺ����X�tv�-7_���}����	� �E��%�ύ����
G�����HX�'T�_���b29I1g�LR��
i�bj��5�GKfB��wQ�8���M�U� ����Bi� 81��{��Ř:.3S־`��5yw�MIoc���͊t��@ ��2Qo�K�#�3�P׏�$$<�.��1�� �dt���e��]ji��]�䤤�AA�)eMV�cS�G+�]���F����o�J�Ej�j^ơ��	�ABFF+ bC�و���cd����c`�YuE�rE�$^���x���8�.��o�������Çr�ea/�\�#Ƀ���RRݭ�d<�����X?WV̂BC�J3�.�� S}�����xx�y߅����xR�"|�{*v�E�6����N2��dM�$ "����:��u��p�'���1��Y���qI�n1�.��h��w]x�L�08aac��jh�ᔊa��߾��?���:5��@1;m�i������.���"Ǵ���v؟)wwwS3�UT�lX�"=P>/��������?,�0{�T�Pb���2Ƒ��O�\���ѱd����bQ����
)�������[���$�܉�sFRR^_�G9�L���P�U�����3׏����h}���pBt%-��;{{�1�p�בP͂�4�����H����& ��Ķ�@����丸ۀn�X�;`�4��b��7�XD$AUD�p�x�M�XՅ����9�<�a	"��A'��ǁ<r��}?5-MlӶ���X�����-��u�;�`��_����؁�gUh�P��3]6.�\��R��j5lF~���5��z,��W|�a� ��߿���F+�-;��8����^���l6�P�|�S���o���ȏ�)Ojv�0�Ǿ���R�?�w�(A����i�?�C�ʪ(��kB��<Q�����x���͛l����6���Hx�c��ꬼ���#��y�U:+��d�F���o����&��7�U��{�Y��Z���K@Z$3��l�f*Э�2캿%��a`�C��45�Q(����ƽi
"�q_ޕ�͊�ꀽ`��.������2O��m,�;�S�V���uB&�/�rr��Vb�� >~���]?M�� rwqa/ 0,l�wL�C������\��Ύ=�3B�{R�|zȱ�/��2y8���մ�	��ǏHV�¦��3 ����kH�ap�)����������M��#/�Ў�! #T�?;_+�?�lD�l�ϟ�Z��W�p��'� ���a]�K浹i�j�!zQ��
֛Ӑ&�_��ؿ�玦]��WLj`z�`��G�R�񉈒�x*R�Ӄ"�># �ɑ��	��M���g�n,�.Όc���wE����'e�)����W��d(��b�z�}��(���*\WG˅}��¥#��ޡ�DEC�c�o&d�f�p�<ic�-�H��GD�e�JK�
�Ջ��*�X��r��x�?%��A��q����X��4@A�_7�x����F5�>����j��zoo���M<��0�ѡ�4a���s�;� ��TE�s�~�%gF����嫕�9�W�)E�>m5a�� �Z�?�͞q��ox��w�޾��Tm�E�����2@4����򛛙�N?���Ȣ>���ߦxF49'���g�W���,��z|����܍�^���D�ʂ�A�}şLsFMC���������D�ɩ�?���OR7/a���n��w~JNSQ�ӛ������$3�XTto����ӌ "Y�Mi��a[�H�r�A���9?"����cz]�()���8�{��P�?#8�.]��|�-:���qI�a�W�����x �_%m!Ԋo���<�7>r���=�`1j���ʳg3ݨ+�| m�h����=�x�+�X�0=͑X�~m$�y�n�A�׸)V����ak?���HF���R�80�v�Z@�׻���v���J,Ǚ+�T"�	����E^��&� �x�Q[AA��桎��A[=��4@��W&�-�-�sssw���ц�o����\Y��(��9��ɓ��-lШ;]����I�z�Q�f�v+Øm w�mR�nx�2\�%%��͝��x���(�ϛ��5����v80�J!���c S���Zf�	N�z�o��ō Fi0��5m|i1w�0���dX��;���ɢ�}��S���D�1@�����Ǔ�?����,U���ٳ�!�;Ċo�Śv�2��EXh��"� ����;���zZ1_`#�;�Gϗ���}��x4 XZ��	x���50ͤB젍�?���-l�;�|Ά�z��Q��C���h}IK����8�q� @���FHXq�^��t$�oٺ�z�ϐ��I� �e�6q�<��<�jg�'O>.];/ݩ�XA�֪jw�{=��5�l�*�?C�,��C�p-@Q�5������~<���Viԋ�r�v��K4r1|�Xh�s{��CZf� �8"�_���@?T��˱
M�L�$���&֔�������rv� ��,`�9�Z(�®Uoq�����H���}�_5���pa+���gAE"L�LHL��7M�w��"kG\���g�b�v�,ZH��o6�5@}�Ν3������������A� A�͆Ã�/���K6Ӭ�QSSϣP���f�wx��[O�W�Qȑ ���S�����Eg�]��H��ڏv�WM���=KSRvu���_�3֟��Nت��$�:2�p�.�!��o��tc,�[����"6�p������E.��P�\<�k���s�nIś��P1I�
��}ĊƂ� P@��f�Z��.�&����*	 � �y�=��Sc= -����@��w�e�ͳ��4����&ѥ+W�AL�(_R�﯀aH�>��GeT���Ӣ���x'�qR����MN��f��C��Yn��ː���:9�����z��y' 0��zV�^7�:���%ߙ^)�Cj�w�9���c�v�sk��s��WU�C.R_<���7.?L��{u5�'�}{nD���g�rox)x��������P�7�5�djk�~��Iք���܁K~b�����I�ϛ��5πL�88>:6��@��DW� 8�&9��)z�DFOHx8=U�I~*GgqQ�����p��������~��תh���ϟ���d��m
00���)ukcP���#""޾��^#&!�WV���J���?>i�v!�}����njC:f�0�M����l�z_2��`�^��O7��a���+������E�Bq��Q��Es�\�~ah�Zbb�ij���r�S>�wgިE���TU��H�5/�L�p�>qr����^��f���3Ʒ0j�T����\ķ\@���п$��x����Pa3�k���.�;��^�}Q�@Q����%��˭=$$^yyl�UM8��[[q��8R!�Z'޾{w��=/�ѫ��'���kS�l⩩�=�.LHx��.vW@@K�@km��OM�f)�98��KW+�pv��3��H���ҏ�����U@�r�22.�Lw��� �e�狃z��O������llO%+b"���,�#JQ�mX�E�:��[�O;%�	ܥ2+D�F��4ܡ���|�3t1>܎G�P�L}w ����RTB"��&De�$3d�U��{&�J6e����&+d���#{޶�u����������~_�9��z��\�,mx{�zr��IA��!K�u�ۣ���I<ve�b%@o~��b8���0U_O��֠�`΀�`���ܚm�袺u���~�N�c���e�w��Jv��m�(=�7���;_�(G4g��h'�n�V�glԹ������=|5�;u�}7����ݰ�[��$�������L	��E�gT����d���77-#���坍��la�Gu��>{�qNAY9����ˏ�1E����ca��g^l	6L�Q�U�R�k�~�/}h���a_iPFj�&P:zܟ~W=�ބlO�l}專����tA����S�UTZ�хy떐���O��)�1����F��!11)�8��\ g�͛7�R�D��n�����k�����k �)?9|�Ǚ��n^
�`F&��X� �8i��Ű�	��ImH=N�k���d�Nn��, or�U�p���c5㝺�-K�TuL�dqQ�T�'�\�MW��Jr�~�I�Am5$������#�_/M������Wn��pS��>\�GL=��
_Sȷ_S3��`� ^�P_@!U�'�~�$�$H0�{(�K�.��9��/|���XY�Ӭ�Od(fr>��Z\S����E[[[���N`	�!9��ĵ����)2��.�1<U\�ǚD�i�0_�f��*�r-�ͷx^J�}�쟟��C��nWCn4��(+WPL���5)
�ݥ�3�$#!Q�=�ϞV��BϽ�N������Km�\�S(�<<l��oD�pTUU��ݹ����,Q��x [~XDlG
	�%J��'X��sx_���l��̸�����1M���mk�~f**a�e#����%=z�Ʀ�����bi�E�4���j�Yj��]J�M�,--5�:�y���J���e�������U�e.ґ�?-����F�)(��x�ot�Q��:��IEE
�{��b�3m.i��%eW<[=`�x9-ap�K�	Pkتh��(�-�VZ,f$28��0�u��p�[�pӰ6<�.J}i��}��;zRo�<�i�c����j�Fg���_��G	Ga�0$W E���5i\tᢘ��&�z�ϟt/sKG�,+�)&��xx^ھ:����Z���?Uf-���u�F�
 �b��~���C66E�X�������M}��3226��NP|��"5� U�n��2h�9��^m]92�;��  ���2s]��HN\�Wuc�63��䖌z��\��ess�xb<<o����]:�6��6�Q�*R�ih`Ç����a��!���릋4JJ�&.�J�S�u�X\�ɽ00H�5�Ǐ�}�i����y��ǹ�ۘ�m�=s��
����!ûuM�mOq��Q������[�d;_����D"S,ioAKY��F������R]��q�zò"<�b��OOGƔ��_�e!L�ˤfc��dT�u�k��~���
���mX�&#�lH��	u�f9�z�\�j8���|=��y�|秈K�"�?�O� #)!�څ2�.�!aQVrp�b.A�1̣�Ly�N�}���@?����s8	��߬�<��	t��-V�A �xx�����֙�K�iָr�y�6E/��^!b���hg{{ʒ�{���g"�|7������33#G��
R�3� BF�`�b':`7��K��s�\s�X��?�-dj�Է��j�9BD7��ld�?�6HGGG��dA�	7��+�r��OF 01�bww���J/)vtL�����b����`��/\���
篫���>d��vwC��.e��cʻf�5n�6�7ǂ��@�f��ճ�_����h�j2jʮ�� ֶ��7���+w�>7?/ޮd�1Q-�c��uee07>3r�/����t��%^+(P�md��m|�ae�0�K+lE������7���������/�.&�ԇP���2v����`�"w�������#�b�p�3L�NM鼊�T���ĭ�����d:�����O��4�I���/S]t�..)���UU��{���!\����U�WK�F�
�����b\�1������3ӄx�w,,����"Pbc:b#"�y�?�IH���f�n�'�����N��1�L��i^J�loP��Ź��S���~|vx.*@����RхOw��`���mz5f��J�8e����s6�1.Yn�H��u_JJ*�]���+�����dL��TX��#��ts]سe�^��_�>�''�,�7 �����Y�}}o�F����{�y}�UyNF�:aGHB"��M�j�SQQa���
k 23�78�1oߞ��nq�=�L����֤\�}țk�l�c��x�ztt�<���?I��ʈ+��u�D��Ru���D<%
�#*��)]�wv�f���$��>���Mo�����u���n���Y���?6���Y�R)G��ir�QO�e�
������<�n�
8�S:^�X����7�@���#�R��Y�ȹ���q�c6�BBE��������HIք���]5�>�ܵ�~�d��� �h��Ͽ5������+����ޥ�>=�{���`�f���B���ϟ?��f�o�m��o"*��'��f9�l�FGż�Xh�R+�;�mgHnEe����' z�.�o�܇�j�yLJ'��#ަD��aҭts,6���t�}�����>��[ ��331\��M�)��ż��5�����C�ax�x�\LI~/HK�:@(���1%�z��l%�o9\����ï�~:')#C���UQ�&�ǩ���gNN�L�N�Zw�	�& �_� Ac�^T���#�����U(&��G���>�j�m��i�$K$/��Y�W?�5u������Zļ��7o(����G=O��x)�u<ksQ�����c�3��xE
����/�e�(���jmm����|EV���XbN�mlRX˘5+�����o�����C&D8��F�m���t�~! ��Ȍט�:���zW�T$'�t|0/�h��$>�����/���N�Nwu�Օc�%~����R�x��]0�@����s��g|<�]���҆ �;_��y9XY�@������*�]J��oYXV6$�4�_�ʑ0����ML�fl�ss���g�������ฅ��!�;�ӄ�N���w����b�ff��o)���?��"�з��6���S��|��K(��?SK�������s�8�#E����T�Zf�f��I�.���H�!�>QlB ���5R��������%������#����ԲO��rNH`��{z(����X�����w ��o���捛+W}Ғ΢�%>w���p�OD��8�����7z��.���LT�;@8��v�V﫽���\L�!�Z��$~��Cv�,��U�/��ㇾ�f/;>�'��YR��n6��4��(��F`�Р�n�J6X�,�b	��Z�!��D�c^Jan�[g30�a�7����d�@a����~��U�>�'�

�3l�#S9�"ǂ���C�]kN�OӋ"���{�6��e�̯�q덮*���2��� +Tjݫ��w{8/�w��\��S���zu۽`����|���1Q��3��{���%$L����5^� ��Cκ:�M�-�hOמ��^��mJaY�W���md]�ʬ`�K�iT��<�bm���/����M=�S_��J����B=\�n��Di������3l�G:�	��_o�j�7=���u����9�����������* ��n�(-�9����Z@5&*ڋ��A@�>΁��F~�՘W�$쉮����܉��wC�2�s�cc��OcZD%3��hQ�����q��z��W�G����/p������>��t�A��hu'#WO��_RP�^2�-�l��}��o�*�� ��Ζ��߰��ܫe��������۝�JY%%*���O �Q�Ȑ��G���kw�O?��ןhȃG�a�,m^`������{����U�[�yo[��]WX�෾n������L�ϗu4WQ!�R��uH����V-4o�玣���f��23���ӌ�0�E�C`�j%����ɮ�7o��8�������=�8ix��FC�h�?�224�&D�צr�_Oϋ�gsw�*�����'x�p�֭P�pDsC�e���}�7�+0�jCg�%�Qo~n�{bbC�P����C��W�q��}Y���;0NE%j�ϝP )&}c�e o~k���g�("/������7n�³Q�u~:y�T�ߞ�ۈ��홏���-w�	�܋p�z���`#���fo��Ȩ�F�B������|������u�'o��u��x�O�H�u:�e'���7H��Z˕���K��(³�"�u�)��J�R���y�󪀐�2�J�N'J�G�,"��#<�j�r�����b�_%��Z<��(�ذ��j�*	{U���x�'-t�pZQ��˧�g�����I�����{�H旟��ޫ'Է�Q��X���=�bT���8wєzgq�-<)����^3��S��	�ttu�ȫ�)��z����潠%%&�ۿ��\��\���k��zJx��ϟ�Q�Z&V* ������k����'lR�I1�@|����*b�>�����y�ݿ���4����5��W^�^�+�%����e
�cA{w,X�1�W��6x����C�""��j�cx�?w��d�g�6C�C�WKF[9	��Z �[�����@&�P`�D�U��t���-G F����F6i�z�%�����a%�b�6�&
���Ӊ���-��GF�l��������11E��=��<��hSJ^��HF�
��N�r�0q��OTTT:=�/�
��9�wvR� �)(x
ܰ*�I�@x�-;%�::6ix���p��E'z���E���7���]-�,D�l�P;��E$�g^��ػ޾��㻙99����k��vu��l,T��,���ݧ�fӑ��v)8�QVޫ��ۑ-�P\s�P���/�|]��~)��J�F����/�.����4�rS�rxJ���aQ1�ay���H�	|T@����^6-b�T�D�1�}l���EʓGO���;m�cm�D�j����F��yX�(f����N���	u�UʌB|��å-�vh���ba��י��j����9��Y����K+@�IV}�|uU��@|���&W����j#x�I�����g�u�:)!y��H!��55r�c�A(xc"b�i�ro������V�?��x,�wԔ���k��O�Kk����:D�^U8I�p��⧏u2l���p�a��j�DDB�������}I�	ВF�Dw[�������f2x��:�j��&���N�4-�`�@	�>����+���N�)B���i�&��j!��0�ћ>������acb�49{��]W��ח�͉��OS��bg,���vT��IJI�����������>���'p��A��1T�S�SrU�;||J��8����՗p��\{��i�t8�
`��4�w�!�^o$N��j
+��_������7�"���nt=�sr��1~�:��,%%��ȗ�l�zO��h�qqq��y���& ��2w�ū�W�L�V@���a񤵮��p������K���z-���-�K���~��Z�������$@�)�Z(�dU���.��nFU#�J�|�#J����-�Z[;���9�j�{�6;�Y{�I@0:�t���'�DA���'���ƾU�ʷڭ�5��p"�����U��F���ǥ��c�!"zT�Hq�5p��k���'�k:�/޿�����I۝f���&��3����!\R� ^v�Vs������Up���'�
֦���--�[��X���.������W'���<N��V�G�4ǣ�)�j��"�
of��8��!
��#k�H�A3G��?Na4R�R1�Ϝd���p�.���o:f��$T�o��Ɂ3Qc1�O�yG�SX���3$��N5���@�}��㶻�LeBL�+�l��;%��@l^y��y�����o�{t����;K6S��҃)�߱oܴLM�����\\��>�� ߓ����ڪ�v����d���څ���kM^��F.�f���e�KJf`�:�I���5�Ç���$Й�x,[)3�����hs��$�ū����X��l �q|!�ޝ�g�<�Y�x���l?:�����J|�����<�g/�P(�t���໹{v���}�{�	,��':����a:F��h��K�)��:,��V.q;��/gP�	�P�(l�x���y0O��ܠ��]��j�9����Ҕ��:�F*(*N�՗+���j��[��I����~�|���s�٫^h%���ӏ��Tѻ��xI���&_ji�J�q�GYtW��Ƭ�]:P��<���~f�-L��JQV����x)x~��EY���^�ќ]:�w��S,'g7�ڧҪ�n���\�s�m���I�h��])GÏI�dJR�(4oĕ��RR��@"4nͶ|��a�E��	�փ�|�������LCC&'S��mh�s���N�����r�+�����q��]\�|�i���U|��Q��w\/�_;?����^o~@�)��%��r@d�Z�R���A�+�oX�#�X���H!C��YQ�f�A\�6/%���444tt��C !����>3���;�M��o[�����Lťk*�b 1Qh�Q"��;::��MS3.o!������+�-���[`Q� ��-���s9�z� 1�����R̗s��$�c`���]1�m����9=F��"��{��������}D_w��J�55�DC�_�F�jO�-��cAs��۷R�1q Xo�ӊ�3w�oO644��:)�)�����P3�������#Œß8Q��龗�==������	a�Y�����l��=��Dmx�v��d
] �Z��B����ş+�Wr*�
U��{'�2Y��' �����K���&22��g]UN;�����(0�8�:s��3�����́sa2ދW�s����{י���l��ū��&Cu+�
��"�ACG�UV�� e1�%))	,�榥��������o �����`S��R��<��� b�13#CB%��? �#[�v���N��kx��e=zz��ǹ����d-Y˗/���{r2���~�K�!+յ��-1 +ˬfY��*$����:�9� �8��55��9
>#
JQQ��9Ccc!�{��l�jjj0��n���n�A}���1��MllQ�������mo��;Y<��jF8=p
������+ \�	Ÿ�6��B�oe�m�G^��9��>��uW42�B���@��|�Ȏ���q量�&�F��-�� X#v0�o=n.�%$�a��0Ĭ+_і��2/�����t�kc}]�ͭzs�+�ˆ��{�� 2�����376~qF�x9�����H|(�!a�� ��db8A4FkiBTTڑ��G�͢��r�?�*"6�3�����F!�� h��F@l�E5��X����v^}���%�%p^��_�	����� ���˃LC��y��K��z��	�eV������f�����g�z��Byt,lؔ�W�O�^�]z\��q �^��{9�,�g�6x��ʢ�A��|�=�����zsQ�+.*���q���l��b�7j�-��@��Iy��d�`I0�Ϥ�=�E���\Xl=}���,Ѓ��)(w��x����T����(,���*7�E"筗�<O-�lfj�J���{���'�h�-�dK����6�|���m?41��9��Z�&�����'rq����Q��ˣ�{�OJG�J��,z?��M~�݉)�L�x}�g]&&&}�FB h!�}��t��������'�Z�� ��@�7��uq�����! �4�-����W��Y��I����ii1z��N��I��5l��@lhi���M^��u�JYEEj���E��=%����+**6A�n}�%�,�]�`<�~lF���Sa'N���	��խ:�������~ \ʒ�����b�kj�a��"�	,cz���H�����/"$0��t� s���CmcL�=�n���Ds��!	l:�tl��A�u�x��p�isT�.�t�r��G�RVa��	��O���e�33��{G{��]�/�҈?��F�o``��}��,�636�/�7������CC���lL��
Z}����]𫫫)$���d��Ʃ��6�	�8>�J����c�1����I�k^��u//��J�c~^�߿ƺ�x&�2��̀�����h�Z"_����ʉ*k9���y(l�������Aڣ�x�x�no�x�d�+}}j�x^��O�z4��H�vvl�;R���g{�N���MO�{5�<%
T)6�ǈ\UV�i�&S��xu8��D������amTE�|<<�*��~G.s� [.u��jseJ�Z�f�%7�.o�guٔk\P�ţҚ�m<���x��X��$�,�vw߁'��	�4�8���*�O�(A>�f��w��ϷuU�z��@ZX0�u�	3��]yY�c��O��J���W��z v�����~��(ld������ p��ٸ�V��Ǔ珋?�˧:�i�4CEEu\/_�엗�/���U"�u�qe0��E:���-qaQ���;0�3P��p�Ľ�=���r�p��ߝ�����h��+C�Q���.�{l��b��II�r���Y�}2�Ta���XWxd$�e��Q4�C�<���H0X�O�j_�@�	Nhʧ-
�(�������)S�[��	��$e�Y�m��>���㴺
Tf\5 ���5B��-�j?ss��A [�K�7^�؀ڤ$��V�p���c�u8�]���xi�����.�/� 2�3#��ކ�m��[	Ę�!Ll���X�6�&��@�,��5�2����#4�o��ҳ���:M�Ƙ;����e^��.h�P����:�QQ%^(�Mǜ�6L]]]@��}k���_��k�����8��%��p�"�FB�Zż��}������d�\ �>1�����Tg�[MS��-�6�H#�������_�_b)q�u}�е��Ɛ��l��,�^ݸ�k��c(�0�~��#`��ջ����M��8<c�/-*�3�,&�:��V�O��O7ס�P �B�?&i]����Ba����F��.P�F[3MYP[�A&W�6lU��$�^�̐ŵ�ɚ�V��->gk/���V�^�����ⶶ���?������[�ÒÝ�X,�x�}��~v�1����@�\������tZV6aש.l��K�io�v�>�e#����	P.Rϔ�ը͞����)���n-�D7�����^6�f?�p+��N��[�`�5�1q�|r���N���Al�V���aE�4�K���,m� �v ������������ݗG���� �x��m�"M/�-t�z���'4�奤d����H@o˷~h �h�n�$�sV0~P__�Rb��"��,%�{{i�qŅ��)e��@��Ra�n���7���R�b�_��d�6��u���b�6����l�hx�����"1�_���z��)ҟ]��� �n��yj�@�$''����y�}���3^YZ��f�w�oĽ���� 6(,�o����~�	�{R��}�`�k��RŸ��D��3i��Ħ~"�+R��1c����ޝ1IYY��鿲�����1Q��{�"T���f���|�Tđ���*,�ޚu]���>P<l�������Kp���u�ن"����9X
����Eaa<�piˍ�5���k�q�M��* ���1111A9�^���R�uk,�ek�.�P�˅u�r_�M�c�N�t\RZ�hcF�2�i��1pU��~�k�ݚ��c�3�jU1WS�2�qJ�Υ�zx'dCMMms�m� ��ݳ���e���.N殢��b�*<�k�!�q�!���_�	�\�Z�0;�}����L�����T��F�؟jK���`��z�R~>:2::q��@Dg��-`�T+�����랼�>�ʦ��Oxi�amCC���S��e����c]���),�k.��*g�/P������)D�<z�V�jno464���N'�"�6<Ώ��X�8����i#����"����///׃�O�IH�5�L���Y��=w���x�<�j緜z_d�7u|�nӼ���N���e�StYZZ��D���[l�{JN'6�cq��)&_�[f���q,�5���и�����\#EEE�?_C=`�(4$<��}?A~}�7�y/Pummmgn��yy����*�(ie��}�i�xzU�Ɩ����W4����`�Rx��躑���ܚ�G�An�|�/w,�Za��~2Kv���S��yxD�t~),P�G��7Gz%U5�����i2s󜙷ɢ^�H�;�� ���Q6~��imf&&�l�b�aU��
PS�oR�C���KG���s*E��|\���}�$#�[DDJYH�2�����-�M��>�$e���J�_\܉N����:h�#I�C=W���+�zmK��L|x���%3�����o���o�̚��ܘ�U{h����w(��Ȩ^�}�UXЍ�Z��oz�M%�W���X
���`A �8��� ���{��P�L��jCVv�ߏ�|s ����[�n�NNN�d"h� ,N��O�I]7��ݻ��x���$p�IH������$�'E
�;��cPP���럱�t*��o����6���\@3}L�:Ě���b�U5l���t���&��"�sA%�}q�v����r�cL'?���?��34$���ݸ�V{���U~w��i��A��eG -��Jղg�h7W�Ϗ2�OD����M�+�!'=Ύkω���2��a
"��<������(�=##0]��w�ebf�oh���LJV^�Y�sn,������vl�I����4�����5::�2��o�6S��cFc6f*e���� ��셮a�Ê��q�^w<���<�+�M�#�v�B�f%��vR�6�;LF��8p��ۊ�9��:�S�Zj��w4�}W����v�:�u� ����dg�0���%�1�NŘ[Q���"S�qhS/4�<;�=r�)���J����l���V|�Ǐ����211��$+�CDD$r�M��YZ[�ɐ�� �D�@����ZR��tY��~����ëҀ�>���461��e���?�0KXW�����/����=�5�S�yx�
{�]U՘�Ö�������H)V5<���1g�q�yL���Za���Du4��W�<�Q�
�<�h21�{>�̬J|�q(EK��v�nw�/$2�0�&����6n;O_�*X�۶�8y�e���t�_������Th��c�]3Ě=d*�J�wHHJZ5br�h��o(�o���l�Q��+	�d��LM�$��TL�e.]����f���XVq���%�N��El��R�㜧�f[��(��===�����,~���~�/�-M��4UhԔH�d�+�gJOO����0�'��&�m$�����1����ȥ����tFᤈ�5@��f������CBC?���ږsp��}f�À���\Gɳ�i�\�G�ڹX➓E˗���&#��>�塥���0QSV&������TvΠ�o�����������"nǼ��o�v���f�w��j �����(�y����i+�b�u����aw�Ȃ~����BI5��������y��w�m�"XȞ��,���/|6������RD�<<jg�������߿������3«��[aI�����mmYuX�p�߿���8M�����=4�����k�VWW/���tw�/t܇�ȩ�o��Y�����j�D@S F��&������)�^d������h���\�ɲ��������x�ˤ�F�1q���7�P!���/_��Р�˟��.+p@���\l�n��q5t%���X}����R�'�]	�p�z4
.F|����ܛA����'@`��>���-dq ����ӗffLD���(X9.k��\7����h󻵡��D�ll�m��Cո	�%�D' ^e�?;�����8��]X�CVV��c{�r�z������-�%7�� 0�͸<�����#e�}��F�!@��������F����Pݬ|�L���=96:����'�D$$r+�B��wQ
N�m�G̬�.����$�`�]�Wsv |�ϐ�'"7=���(��K�OضO�#��8�UL�:VÂ�nhh8,�wG`E��[���)mh�p_�]�&)11����ܣݣ�<��zϮT�VX3�qV�ౕY���}�D���LV?��o����^�?d5'�ϡ��V�d�/��F�U��D敫f=,�x�Db���<��E��d�����8ԉ�eK�֓��ʘ�N�m�	X�e1��-v�9��<�s�:?�|�t�Y�pO�3�\ ���lC��p{�q�ۻ�zt�Օ�b5&8Ь��/���v'#��j��L�ѩ�(,T�e�n*Wם̽}�����(���Y��^j�4�}1?�q ]��us��A���uy�sf�,�E)Ϧ⑍&:��c��.¿�jO���ǀO���so�07��,J \�&k��6���6ȓ��
�Y�i�Y�&��X;��jg��'������(����i	��ӓEiT»/��oKZ��9�M�f�|�*v<T�М�&����޷�muV�>n�z���EK�MOlƕaQ2��)#|���^V�@��6�㚍���p�_��*``D��b��oEm+���I��5��v��p��ҋv�}ظ?���ӆ�n��om��y��v&��f%�Z]]��R'�\��	P�⹘ugm��4�����+�Sz�I8�F�N�mX:�=
8�<� ����$l����6obv����[p��%��]�{�k�p1�Y�%2���qC�Е�,^��׼W�R�#���ݻ�:�R�^����;����Z�R=n*�j�X���D��	�����U8bi�5�]=�;�~~��W8c+Y��#M�5�۬e� =��ބS�9��Ӯ䩘f��`-lN�EFJ����P$B gW����V7��Sa��!`�15�E՞��դ�{�$R��\�w�5��tnN�hmD5�imT�>��t))(gi%@a0��.:!�y>���3\X�CpzT�e4Zb� �֢�O<T��X�K��Dʌ��#X���h�.�
�r���o�L��L��k�#x6��O�2��]o41.�\��&�HCv�`6H��z\�ƾ��a�[\:f-9�0����Ó9��o��l��妥���>׽��k���R��+*p$�FQ`����R�aޘ����ϨwS�(����hPw�S����b�����$Q`�|�1؞}1Q+S�ő�_mF�n&�j�;�J�I�n
��b5�U�u|����N�q}带vW��'�S[dE����r��b6�P�s36�x/�c1�:[����N�&Sq��|
]`ik���!��F��7�� zԼ�	����cocc�5f�Q��;�
���]�bq�M\����L���c4� 4\r�%<�ތV�����ua��ݻYĻ&�q��hH]�_������`-k,�6������=��Nl���x�2��ԓ��bRKL}F�o��οZ�Y�%c��tY��Y��c��#�6*Vr��G���7j`�R~)�l��Q���X�����Z�8�ujv%^���UZ������*�!��4�=�S�d7S/'�5��.˥�l6��ck��=;�u�t����5=\߼I,���OaJ��a�(؀��rv �g$M|"'+r˪ېu��6�p&?t`I��9hb޷J��Sſ�����0U��N�������ѐ���oI��a|����5���?��ø��ۂ� ���Wk��')T-�m,ϲZ����*�#/�w�m��}�PY�8a�'uѢ�W���崄��Vp	��	�58��h��@���t���	��gϞ��Xa�M.=b1�#�_�����'ª� ����[9�.�p�XN"��]f��;�����qs�I��'mK�ȴ�l~t8�%u����9���c��k_��{bv�������v6(�IzG��{���^.I=t`���K)�v�)�.��?�
y�Y����Ό�8�8?����>+���ϲd�v>R}��xc�z�jaW$���*'z���S�t����Q�l�����E\�i}�^�r��X��01�@��!8nᄺ��?����2���ǒ���;3K���_V����S�'�Z�=[��:C���������7�S��|�ˢ��f׉1F�߸86h��lܼ�,��7&������p.R��1�a�L�J��H���ROR�*�y<P��1����!�!��Q4��d������WW���J�+���L0��}9��]â����v:��j'%��X�|�}>-��촇��Q��d�Y�����kठ.ׅg����k� OY����"{=Y���/l�VQ��8[b>^/'j�o<�2a"�I]A�sS��%E����9+�u�>2�����ץ�&=��;��Y_M�o8�Ix�v�i;�Ě���f8��l���l)茎Y��t<������K��2I�ڠ2ȴF���^F�����?P�����i�Qv��r�/tK ���[MO��Īب/Un�mG
jJ_,�O��(�{�w�Y?(�����<��d��v��1���ʽK1h�#=u|�<r�.MWx��������s��̇������{GlA�2�TH��S�t�ߤWr����`�t�܄��䄋m���~m�2kh�	�·���*,��`}Xb"�_?K�8#�X{�7���pCN�)AדY��]c62p�x��"��+�T� ��kN�V-�AY��� B�t�2��ɿ�e3��z�K}f���(�h6�7 *�]�\�vť�Z.��w��]L+�F����ۯ��/׃#�*k�+�GŢ������Z;E��G�%�\�
;c8�|S�8p:�/8��?� YM����Mn�P@�R���>a���MV���u|R+/O���7&+M"���w	�Ty~��,{�հ3:�-
*�_^^�>�Ώ�(��eɾ����x>bH&���-����`.���A�����E�9&�|r�:�d:��Ur`9��XC���j&�ɌH�F|K����/��6�܋�Mޯ�b���E �ʤ^�+���`��������H���I���6��徴�l��\�>4��qs�����i���^���6��Yd�삣�. �����|�f�i �s������\k�ǥ�G{+sp�+c�Үh .�����1���c��"~^������Ͳ>�����+�/F��Cv-�AO��y����3�ܦ�^���B�L�E��n�?y�6�E"En���bz�Ռ0���@8t ��Y�'D���B�g�x���'��j�,�����ؾ�U���œ�2�t3����	�я�b��*����͹c+ٳ���~(�ߍ�U`nI����T�3�wZ�<xT\�\֊�����N��ë*Y�i��7$#K��ͱ5m�
vUhe���>�y�����ut����%#W��?��n�Ц�	߾�Bu�1��3oKg��HA��trR��:�$���Ы��'H���D��� �!�s�i�y�*�ǿ (�&E%�ǩhT9�>Q���H����.�}B���J1ZR��r� r�|��m�ժ&��R�9첡��4�	U2�=SXCН{)�u�{3��3t]�E(��XТb�$��w>����	~��>�f�H����dw��^��Y�C*�OPXl!�(h!$L:�+���ܑ��O�9�o�4 8&����I����{��Փ�v�.����<���s�^�/D�ْQs��{=��[-d�.�'��R��r����� O�m	��C�\���o��>:U������4�����O��8"�[�m����sw8$|��
�$�J�/�%k�-�[,�z1��7�u:��������W�����F�����a!�oR����{��S�?	dpT����3cDR�/��p��uum�7�h0���3��M��H��Q�ON�'�G
�ܐ���0�@��\c�Cb��>`�o-�#�(�ﲓ�Jr����"�J|׹lPI���w�V.��9����'�����.��ow9�})�4�mZ�����]�K��5��!g��-`+_KG�+�/,,�@B�����d���U^�[����&Y��Z =��kn��5>�υ!liE"�0E����z�D�X-lo��]>}whu�f��<{�'����DV)x[B?H� $��Z����I=BR���ɚpIU#1O�4�A(�׽T<�@�p\%�l�����ɽ��/|��|����A��H]V��BO�5�f�꽬 G-h�" ���V:��i��<��M�BXl3�0����:�� A9�1����}��|(�EC4�3�����`x�>���'1�^���j���F�-=���u@޿Q�t��?X ����ws[�d���>9L�\��|�C��fG��2n}�&����j*����\#�K�ŧm/8 <o�F4��4Wӑ��U�[��C��X�dÎ��{�� �w��޳׸���F���(%` ��&��߀.�q�������U��8�z4g/mv�z�dk�l�6��mE=�ac�����RJ����%��Ó!��^g9W��%W�vc�z���O�|����b0����(/��l�r� '�}�ڬp�hg1��n�T+�5�����0J)�c�K��~%2l1Cv��w��q��5&���J磾*>�Ը|�^dɸ����S6�ƀ�1OڴA��+D�����!�y2Ej5�KJ46}H�^J�M��j�j@|&�Y���e�����dv㴺���(̓�b�G������x����o��p>���:O�K�S)�N� ��5L�N�����a��I���;��{!uB��G봁D_�� @��eP����]ӢJ��Kp�\��}'p�z9��у�|����b<js��n�p�Ť/�/X��8�H����a`�u��mP��d����X���?6E�e�q�Xd���� �ƣ���zͺ,��(��$"�e�%TS?LHV%q^�s��A.�޾X�)�N�m��l�L8u�Y�8>1���@b�f���	8��m�'�|8�������&�8�@�
�_��?NP�6Z�2y����K�����.��v�l'E�ѱ�[�\\�k�:�;k�N�>[�w��sz�UkJ�V�0�qph�i�f��e�d_��M�^�@��?M�6�o�V�8�X^^�����*�R���kΦmq�1��Vq�\�끵���r �'X�����d0фHb�
@E�fО����P���/a����@X�H�1����^����qs�u���:ϋ����3,U��ޞ��C�
ʌ���Kԉ�F�.���8�̂�5��ܻ�9����$ ��:���P�������՞�`;_3��4����l�8�t���Kz���oA��[0U��UL���;�{ O�z� ��ۏ��5UL$�b����G�k�����:	u�]��=����f�3��ϫ�-���U�v�t�����G��#LEB�4"s^�(��]�0�yn-/�*( [�>G=�H����߳P�C� Mh'}�t��y�G�x�fX��?
L^�8��YZQ��O�Odbd�k����3�Gs�V?�2��{=��c���O�b����s��K�1����nCV
�m�%4���ǜe2�ߺ�λ���'PK����\�Y����]_��.G�n��f+�B��ޥr�п�o߼I�n�S��rcgi*��\ͬ��������{�P*?�j-��r��������(�u�b��;\�	4$#>�e���ɛ6���k���|k#�z
u�򕼌�r�V��	Sv�\�),���CS�"�����چ�vn���E(C�&>tt�Z�'r%,<�Y�y���L��gS5�g�_Y_e��?(Z�Y[Ȓ,!��Œ�d�.��{fl�E!2B�$�"c�B�A�mF֑���޾���u�uU<�9�����~Ι'5�|^�����X�$_|�;yK|����t*7��c2a�z���@xY/̱�Nn�ߋ�hܼ�F�0,,�����1I{��`�b��l��	lC������JſcMUQ|��AF�g�ɟG��Aё����oAR�9���n�a�ֺ���\"	�W����& ����h,����(��p�p�⴨~Ďꣿc����H)bS��-1�]x�;� j�J����S�ɝ�]l䙢Zi�Ϻ�w§M�}�bit���b�5��d��~�x�z��<b�a}!M��� �!���ٕ�;���W������+�_|6Bp>S���	,�3#�.���D]7���м�����U�d��`�,��%�����TL��Jg�hFJ�d���E��dw}!���ls�0�j�<�Mlz}�����8�&�����	�崶�:�D䞞��?i�m����'n�y2�{�e��j�����{�=Ī���W�"�M�l��7Z�����ܟ���*����L��I'�Nt�+����R�N������];;�#i��4P�4���Z/�*V�=O����E����n�49R�k0�1�D���o����R���"��C'*�;xt�GU01�2O��Ŕ�~�����K9^^^]$_�z���N�o
1����{
ً8pn���X�"1���~��X�w=�7���`��Zb&�ӻаX������t�'������Q�y���|#Qy�{f���[��ÿ�`�VIx��`n��,M��5�j�4�`�t���{yU�U�z��]C=�� eK�����u9�~�� 	{b��5Yڵa{m�)�F("��p��d_����d$��+��י��J�����W$�$#�h�>D	�:[�^y3�o8J��y�3����Pc蛔x-�LGh��];�!Oә���zJs:�
w�dӯ*y=B � `Y��L��o�q>y=O��vN�\D�� ��YX@��L�'��t��.%O�����t� ����"ybm$��f���N�w�=!���h�����빳�yy_�� C�$����H�)�(�2��F����uyy �6�=���=Z8�5��@��&�B�,~1�5�nskQ�
�_�7��R�6�#i��Q%�a�u�o27�-��{ibڷ�&V�Z�Ѐ�6I��U ���N����p�^�ʸ��:��B*��\�2�:d�)�������ۦ�#�����,��oX5i8	�1��+�~��F���?J��%����J�H{����Yθn�z��$ɤӲ,���@����_�Ov9�[��^�K���fN\=ow%�9Eډuu�BA�r��C_�Wj�9inw��;����P���F)���m�@ձ�S R��a����5���Y���9�-�c:;�:�잻�۽�a�c	���y?�׺�WP.
���:)u�Y
Ҕ�F8�Qq��X��/xTw��l�k�󨩿ާb@�J�������1�A�w��P�r��{�(ŭO���;���g���p��!E���pF�'/E ���7	���F�kGƘ=1�lo"V�Tמ?Pu����P2 L�R"��v��a�b|
zQ1��O��<��� WXN��@��t
z��\w��c�k���W[>�ugA�uI��,�����w,̰�)/�!���BD_>_��_�W���vk�����x��-B��f��;�ݝ��F A��<��0�Lj�L{��A2���{�����5���͕������/7���ef&/��}�p�����޲�h����#����W�?q�7���X�7�˳q��p/��4�X��6U8��@�晻�i�G^�^��>o�h�&(��X\O�;@G��?%L#%�����=�X�d���UE��mѦ���š���L�C�����ؿN�(@x������:�+e�(I���<v�)-��m<f����s�C< ~D����=1|1)W�Q<sFE`�#]�qY8�t�~�}[a���ֶ���:Z�O�lw."MA��SSE����ERZ�j�[(�W���3�w��������:6Y�LX �@���B �Ca+m�����W�RZ�*��YXn�;z������镡���Z�[a�������U������7T�t�U����V<-ť%G#����K���	'�����a����NCw��R�֠�P�n |�ꟺD���x�l	��3/B�?���[�p��F�2��W�~�����|u|rD)c"��� Qj�n%�<���֧�Z��gs�� z9��%�O��
X��K͈N�=aK�/���l�l����7d�9a���$��PL����������x�m���������
�aj�5�d WD�+5ˇ���>vC���&��HJ���I���x�s'q��?��-���&c~b�RS{=��>�ԑ�G�yk�J�=E�)��w�&?��.:4}}�𚚐?�p�7p�^��i��"��(|��wv.��'�;y�ޣ�����ȴ�R;�F���UA�i������4I�L�or�(}��E���%��e1���d.Ö�����T�����tb�5�>��卮*�
����i��q�]j������^��p����s��GzZABb�+����H�z�_���IkOt�i�\Z�]0+�LP���'?���y����ެ����1�|;ZV�t���cI��������^1��3�㪝ң�%%�	�{Q4[��c(D)��)�!�^��*�S��7��w�x��׶�:���<�� �o����bw�c5��@�~�������Q��2���M��R��xO�IE�`K�X	��_�?A�ܔ�����*���ǘ���(�_��g��9�P�a�.9E�I��o:���W� �'���i-]).��Q���2���/��nwk�X9�]����_�ނ>��pE����}_�d��b�:���9#���`��$c�����<��l����n���Ũ��[#aU�7/*�T�sV?���b^e�6@�q6Xf�Hg/����ޗ����z:���!�A5sz6tp�����]�5��?������m%�Ш+W~odr��B��U�F��Ș�I�1�����wo�^��z�zBFlc�h!r⛋,�� �,1���\_�e�
�����j�H�5����Va�j���ޘ�M�]W�Y��PCxx���~Ê�̑����w�{�������t��$������|�9�
�-�RV_]�0�o���
��RbM�:Mu�}G����%�>��o�0?RkRsv;FF�FGS��g����5���ya����3��\�3�Y��������x���=\\u�@U�S�?��1<r�\��{�A&�D�ZD��N.��ԀM,,:�cz�����A?���0���7��[7j�{-kloA�\ϓoP��NQ(��-�.��n��v�4�<�����ʪ�ɴ>�
�	j^Z-�]�%���\��r�����+ұbE칽;����A�@ll�CG`�s��e�y�1����I��8`$����53��C�?�����X�j�ʄ�7!C���P�U�-f~ē�;��'Ϡ�6��
�x�q�TG�ĝ[\�����0��9D���ON+���hz�S����V���/�`7��?�1}����[��L��,�91J�g�����S{㰁�V��eիs��� �ir6����y�� �O��E�H�y�C�dΡ�U{t�<���&=,��9�s��Գ�hb;������H���o2���Ig&X���L�R���˗/�|���If�D~�����=!{�2��*a��\5ߞ4 f��)����B,
T$1[Mt]A(`�w�q,� ���d�m��0xP��j��M��+�a����N7�_ˌeț��셝N2Oi�!��dy��JƳ��g��7&Ѕ܉�u(#���l���z�hj��z�"G�8�3�g�v3��C�����p/�*n���X�h���c�n/��� `���c�L0�D����=3�w���X)�����?��7�-T0�-v	���r���[�:�M�Q7a�+e�j[���F�o�}����\ �U�xjYf)ův0���А�h8O��w��o�&�d`N5�D�}�*6E2�����(;i�ج��9��c�|5����+`�d������l��e�H���߲� R�h|���(��U���G{���3<h}�'����U�*`c���:(>����eF��=F���om������[�zT�K�`��0��a�N���k�$�J)� P�LQ�}���V�AŁݰu�6� ���]�D���7n��͟L�c�� ���0�g(�@�=-���YG���A�����Ⱦ�(���!�6���\6;���k3A�+�\WŐ�~U�kea	�t���+{����������(���YG5o�%f���xy2e���F���Q�\'a�Ϟպ�Sq���=" D����>���iy�.FVqA[Rp��:�˺��Tb�8��F.�d�G?:@�-��:e5E��i�?�K>��u��Zz$r�#/D�I1�ԋ���>y���?�������[I�1�[�����:��ұX��D�~��hd�uI!�����B�-�&D~L�ޭדCJ�M����iZT��P��/Jఙm�'�9�w3�����8��K5V"��Nσ���J�]������k�:E>wy=C�P����d;�V����܊��'{������%K��.��3��C�A��Zm�c1�3�ޮuK=�����^�.xw(�����АpW��i�$��1,N0-eC�P= ��V?��]�Zğ�V��\����8x�Y9:v������ 	��BAh���.��D�@�ϵ�w+��7R�v>��NP�{����[��U���t&��_E� ��Qg� ���Fa��������yR������!]��4�3�&$�2�:O���%�0���`�:Q�6���h](V��QA.sE#|c	^�����H��w&gq�P,��ܯ	�FB�k<ƃ3�g�� �؁X)H�e��E���>�L�2�4V��5
mY����c?{SC���[�y�	�]<���{�މ�Q2�`���'�xlx����B<��ܒ�����y� �&�xNx#䵔��V���`��\�T	R��9Rv�>�o�J����%:p���mn�W���]+��ߡ��c�����.������߁�9�,bTh^y��>\�6���d�4~�4un�)�d06�:���_V�x|b�i�tl�o���p�r�nS�f}_�݂�<bG�tK���)�<�>QEc!�����@_��;�C���<)WO�d�T���w�H�u��u{��0
Th��ZO��1LE�WT>=9Z�߁:ȁ�K�J��	LA�������!�;j����)':���	�F��	�
����呌}'<�W�D�`0u�c5:UYG!�l���p?���}K�Ch˔]�~h�e'�k�C�
b\��{`!q��qSo����)8�0���<b�30.,����%���6-U0�lA�{�> `:����� ���{��B ��g�0�梚{Ԋ��Cd��G��k��n.��W��l�c�:Ԧ����Sz��S'1�!F
��AI��T�$���b3s�X��1��@G�?������{հg�HD����}1���fsŻ�'�����T��� �Q��/l��wOXC&Y�u=E�w��iq��6]���:u��ϫ����Ȁz~�%���M��>-uV?5_/���N�M���2��.���x�k�������0؄;w�z+�{�˗O���4q�KF�yޑ��D���ص+k+|��HV1��t�f����z����0grF���qv����|��� /b�c�z�sz�`������r䱧 kK�u�?'���$w�=�:��}�n�E�y���%��4�'�-l���2�����o�0�v��݅����8�f
�
fV�9�lZ�U�
��:�P�< D�d-�z��|C�|@�j�G�٬�2�L�'��^�5��Ӯǋ�j{"�s�r!ch��2m֎k/���6��"�	^��ݚw��O����A����ð�_�_�}�j�u*��-P�?�{K�B7�}����������t�6:E�_.?��C�B�-�� qB�Z9��k��'77����0_�a�,FJ�H��?��M3jN2 q����&��
,�����j���V��k ��njw�����&�)���;t�K�Y��v��c9�+�BK�7W|��w��M���4U�_�I浾��"���i@(Mh[ϱ�;9�B�=�Y�m�P�Ձ���M�|�K?=S�)��.�8�ȷ��>�F�]F�6��/a��/����ӓ?��ʋ�̐�ʑH�ZlA�a3����A[��YZ�؞��ǦBug$��!-:�{��h���R�D=Hq��P�n�P�~�D���c^�����h1��f���r2."��������,�!*C���*4�=����BI��Y��&�W���9-����	����[�ƿ�b����rE��B'Ła/��1O�rT���5�_h�o)�VS}H��<�����9��E�u�9�$�L�S�-2�C<iQB�Fĝ���PH��������=4JL��()ijk'��q�]�.���tT�n��+��� �eP���9.��=�PT�n9��x�%$����7 �Ջ��j��[�죣��A�b�t�G:�os���"�!϶�1�:���"�?�a�o+�e�����:�9����#.�3|̝׼ݶ�3B�J�h��)�B���@��q�O�� _�/�~͵��k�~�%,PL���}m|r�� �T�c�@wL[���oL�4y��~�ε>R��Y�/��&��V�Z#�{	�Ы`��۝@5��&{RkP�Q�y�u�Ef�s뵊G�	��ͮ5UW����n� �n	��er$p��j)M;w�h1s-���6-���TR�Ѓ!-�d��[�4~�?u�~>��x"�S���������=�� �;�̗G�̠U������= N��˝�����y	(@�?�*M1X�������'w�r�LK��p�ӳ�l��r<�P|�>}�?9#�#�a��0�2��\�;-q�Z�#�C��p��CO�&-�@Q�K��Q��$ H����J@�5]�#�����O�-�m�[��S�T�{���P�uI��K�n:�S�Ǐj}�,�j c�æW�1�,_��3O��V�N����`A,��P_�;
����bC��Jy=���S�����%��2P<;�=�.�s��N����!`}�m�)��ݠ?���#��'������]�j豗����8֤�zS���Xn�=5���O�xq�z�4�<Ԧ�j8`�:�$��9V;M6��dy=�S�)����c�J
�fV,�s�,}/+��X/�S�[d-�s�,���s~G�B�:��
��(�<��e:m5�n5�c6g8���1k
��o�.oh`�O�Ί.DI;����Qcm��ש~�z�����1��zJ�oΆ}���S�֗�C�L��5��Pz`�������
:���������:����T����0���6Cυ:�ΌA'�����ד)���Ǐ��Q����'7��>Gȸ
Z�~���FdAUD�KB@�̕�F��U��>,mxB�A��)�c���x����U��Zw�!U(�U6)����CҞ,y�i��Y=8�R?�J�;��Xx��KV�7=��QX���g��s�C�� ���N�KJJB$��*0�9b&gp�I��NS�:�p~��f��-HRa�瑩!�Ѡ�֔9'}���Sz��ɿG.��g�_���������v�7Ξ�ZpFu}?@`�3��N���f�ù.����t��Sÿ;v���-_<�)ܻ_�?��ġ������7Zt��|�ʞ�������<�*�?�w(�>��2I�7�Փ���0���N��XD�������1O����[FG*u"ǹc�j*%k$K�4�YxZ&�����!�aCȧV�%����Ә�΀`�R�pP+o�r��؀�s���L���X�6������<r����ҫ��վ�b�b�)F���0�kl��]��:M�e�6x$���d�ӑ��x!5w�7��ۂ�H�z�u��b��f���F�z2�i���{�pJZ��37��@�U��ߐ��6���$�9��������a�cyO�ـ�-nF��}�Pl+��W��q�PrO����yF�&�	����%��
�0V�c�#��M�xn/ �7+&�W�4�c9X|N5����J��#ܩ�NXNٺ�;�=%Ȣ�鎛����;���z���F�,����tc���9ڬ̼� ��'�*����1龜��.���鲇WX;�R�v���}�2����k�u��}D��~'���}T5�KH��d���sd �?��y8ʼ�vk�D�6��i'}��_�2?xo.�P���A	���2�9Z�u�2��|�5%��b��g]��Z}��v��� A��K���[�LNm�c�jǓӴ1�P�`���,GW����`�K�e�`]Z�>ՙY�=�F�u�)�
$�'���_I�����\�[��s�%|�s�@�&���%�j�(�D�����*|7?��qF5����dL�]�>��@t�ǍYl���L~=��[D�;ۣj�{ʗo�;݋��P�EsC��������b2���sA��4�H���Y���X�x]` �B��X���$�$����w��"^��l���:��>bS� ����<���K�"� ���6��LkN.��������*�ث��a2wM��M�	Z���(#���|�w��e���ܣ���}8Λ��
N�l5�<���f�F��c(��O�Si��fP�O�h< {��̞3�C����pyyٓ�h(�-ȱ��E�E�z�\
��j��,E�*�r4�J���`��_opo�h���#.�W��?������Z)��*�R')���&�k�����`�׉5٘��خh�뚅z�����q6��:�9���W��#7X%X����j��xs�V��ሹ՚����u��YVÑ�B�#��3C��ؽ������\'|�f��0��L�m	��	�=R�� ��1���Ǭ�r
���5��S�z]ѽ���r(�Ml��"+ە�����"vM��	h���p���8���N��҅�;/_�����Bp���N�֧k�B0h��:������*k{�����z�BrOzD��}Mcr_�ϱ�
�c�S����nZ�c�Nh��9sT�D�غ�E��pJj*�gA0��OO�49��ߩ�w��i�Й������5�dz� �=�NGze���f!�����Q�k������������-4mG>v�R���qD��黥��]\������nG�`����e�+Va���^�	�j1��Na�T������#�, ��TV���a]-���@�a�}{��7�5ȳ��� 5 �oL�1���z˽��^���eQ�ŐT�w���Fem��|�ZO4��ÇWV%/7�R&�	�khh �FLT��.�$����:����2�+� {9��zpM�dLqW�3�Gvt��c�Cl�}q�R�du,Џ4^���|j�5�Q��X'��g�HZ>	Q���ή�_uH��#�M���n>�0�(Sz�M~0���j��Y��P��<ŉB.��~����U��=3��}��<�pv��+μ�R��<��1MN�R�]=S{��EX��1x_���R\{�[eǌ���yL��<M,؊��P�5�z�H�	�m�E��rO��$2���js���2ܰ�0\,O��q���1��ܮ��������r�K�������:�+�W/�?�WW�`0nh/��E�F#�MJ�[ڷ�Z�;��t!r�W/jg�rqvb9#&�A�}��W���o]9��6Ab�,Kw���km��rrV�m�y�hf_E���ȉr����Ğ�����I��,�}��1J$l���Y���o?�-�������m�����a�6h��\�]�l�� 1��թ΢H��mU�������?��/�o���MRr/�b�X�m��;m\�y��^����>'�}>�#.�<��P ΧzlD!!��f��Ȼ�3�6au��HP,��:���sA?;C���(�;(>jx[2+�y�n�~���ѐ�*��+(�L���^�E$m�Qx�5α깧�R�/e3��[���m5Ǖ<դ�Uᴂ�^!�u�e0	(��G.����J��|�D�}�5r�ig��.bѴ�7/tҴnu��QB(�ڜ����p��o}-H�y�(<'�)�.1x��6Mv�)�޹Ug�k�e_��s�(�s]m�G� t�K�+�K���R���/��4��UiQ<�g�^����{b�a䔄���;+�6M��x�~ơ�=�x�}��,��,����;Xv�c�wr%��I�E}1F��ȲU�[se��>-'�����tY���흛m���������|�ͷ]���&����QK�ȴ9�C��<t���|76H5/5{נ����6��saZ���99X�V���ǘ�e�[`|�CY�tag1-c�mL�~
���|-�����.������ɩ��͇YJ�ta�!�
b�v��vنs��G�uE��|�;��/�&�ԝ�\on���Y酝j��۱Wk�]�]�%l���.��v�7x��B؂��W��r��k��<ى���+���Q������iՙ�Xv��L�	�Mۭi�zQ�S@~�[͜3�-](�Հ/�|7��N+��\%��ٞ
ެ]�8����K	j���6\�b����W�S�hVP4�o��Rl��b�ȷ%&h�%�ViD�iR�~���@��&��=D�}�}A]l5���VO{l�G�n'[гT a��Ŝ<&�e*�"�IC. ��TR��^�M@�=m�b�fA���j��v�-:�8���?���p2J���\���"7ps�e����Xn|�#,;���Js`��t�L�jF%��{�@6�̮� ���䐛��j��"M0SC��莳YE�Tg�4���N�.Hi	1�B.T�bI�����؆�p���vg��J��Ό�PE�/� ��R�-U�m�6Z�m��m`GB+�5���B߉4
'�l�p<_��v@Y��,7����/N��{��7�j��.(�k2��Ȟ�'��}E�w�g�|�ϥ�U�J��#�`Z����z�.���ݫ�'�5��zT����Yw��á����w)�|�oBC|�����K(��/�-CR�2[����������R�h���2�cQʠB��Jd����������=F�bvp������j"y����d���*|���lmU �N�ۣ�����ׯJ�N����ő�7l�!�ב e�g)�)D�n/�!�J��䛮�?y`/��S䖀��Ö�Z?��^���h�S��9��lb��v�����x���H;��k���3� ��`tr.S�׵rB6�m>��J�G%��H��TpH�0�����,t0��%��������u�����Ň) B �p��5<�ۥj;���!�b'!\agbazx���]��\D�zj��{<ǇpǗwI�N�oM=ݰ��Zya��/ª�ޠ�~^����sh$Q(d�+P�řr�I���[=z׏
Sj�]lPh�m��ױ�Ǭ�Qڧ�L:U��,�8[�n7y��_d[�`�X{.ޏ�^��o(u�o�`�fQ�,�&A�Qn&�=NZ�f*�.�u�$.�}aϖ� J���2�\K/rg�%E�}:�X�S�jU��/���;e.�}}�m������6r�#ee���}S�~j}�s�mwJ�=���nx1f���B��ڋG�e���N�ю�}�^�-%���:�˟��~�!���>��&�,a ~>���f��F�+������.sZ��'���v�^h0�e��0T�6�������O��� I5J��|}`p.U��jb��≵���[P��� dk�b���R9�c������.7���v������$$���|__�^�;��
@�"WVN�$w�*�_��fu���!��t�|O�y�Zp��:EԆ�"���j�:�����go��"����\���Td��I�=���������)�-%�/_�����+앒���g�� �8_]Zq��7�k��]�fyR�C��nL���k���]�־�I#��J���y 1��s�Vc��2g��lJ&�����fS�2�h��E�a�4Y���>�dD�-�dec�G9V��L|~���f9�jTdO�'qlP,dse۝U����_��3�[S�@������ ���CP��*��K;z
���W����{����{��]ȝ}Pt��ڂU����ƀ�a��C�d(n�*�Ff︷��v1���}��%�0=�ߦb�#U��"�Z 3K�}��Q�*O�;�����r�2�XYY�dd������Ϭ0p�=K�μӗh>� �m����ykX�V.���^|W��wª�B@�7J����L��b�6��P�3�ϊ�(h�iɁ)����>SiZ5���y(bh+ƀ���M� �A��d7���lz�X�>��rn&��ۀ-(�BH�ٻ[߼��(n�������	0iX�d����[|N�Btŭh��������wte�9�=:J�і����X�%���R�����+�O����Ys�$���| ��~fO����l�M':-�_��=6�)/����ּ_C4@���C����^Ԕ?��ػ%�S��8z�#���x{k���-��1�3�,�gz@��5?���z���髠�`��L�ЁUĶ�?�zH��j��֌���㡊{���[ʟ�ź����F�ܔ�Z�- P9�(Ѩ�3�qZ�o޷ƓK5���(�����V/�DM�;V��IY ��7�G��`�o�M�v�2t���>@�{c��k� ��ŭ���t1�ij�s�N+b��bN�����o��N�
kf�$�b��uP�0�q���d��&ec��������ȴ����:��7w�Q�P���
aP�.G�k~^��/��d5����mC��
��YLLv���R,�^�T�E���z��O�1fAbª�\��_�RY ��2sL��#�6�l=��S���I��+	�"J�XJ�ӝ�����eW���g�(����/���=�X�3,7��ڴ��5l�ak���T]i�po#5��-z�Y"�ˍ=<�u��;��فv$�{"��w���\���Q�P�ٰ��- �M8�c��j�]6���2��~,��1�һ��ͺ���h"Z�W�����.£	'�f��G��Ɂ������~�>@Y,�f����M=�<��?��Z��� �_��0%�"Hx!��9Mo&؉���~�	&nU*������ZTL�x��^���� �ǪfaS�G
_q�!��;��\��f�z�ƯX���&�j�ݿ7�	���
�J�"�������Ku7��������	�x�N|���S!��G����/3C//�����U�O �k����sb�7��OY{ ����;�ϓz�:>�T����GS�!{Yhk*or�]��վѺ0\��y�(ۻ��(_V��F��M�G���C�����LOB�mA���:a�(�V�?��Ò�e?n�z��)!zpʬ�����}�.��C�#Xŀ*�x4�-3&y�����FB�~��gf
w���ͷ��z؍3I�B�c�!w(�k��yϞ�~ u��UE�@w����_k����;r��acph��9(C��ޏ;�76Ԥ�����C��-�33"vF
|k�q�'/͍�{��o�ʣ��`�e���I�dL����a=������A�Jȝ�����qRU0�"}uu��y!�sur��`b����*]H�R#���\c��I66�H�[��#_ۏ8�9,Ou.���鳀@�4p]𖃮ށL��=۠0��s���_��(����K����y�%i�C�2��7���В��׷���,��V�A!��W,���@��t�`s9����%n	 �3��T�D�)O�1L���7��E�?����,��{��$~�7M��6E�d	��ρ��^�����3���ȵ������I�B��0̣"�X�B\���䍍jt��$t��`�7`0Py]Z���H���QȍD�P��c��V5��WH�g�Z#O1�&2���|X�CG�RM��nJn
�#�_����x���>�v��xA��1���ѽ?`��Yy�t��F$_��B]t�UI_Y:�f#w_X���5�m�䏸RU���@)=S���N�I��T8_f�wWb>�HL��j�[��*��A�B�y@�,m=8K#r6F��E' S�V:�3�q�i�|�'���������j,:� n^C�� hF�.M3�}D>���]/S����e صeCB�2H��i'I�z?������6i��Ρc�:}!���ΡS��'��HIEI��F4f�Y/�5�YO�2؊U�x�DH�U���/�s�lG�K�Y�w�1���,U��&�Ӱ��S���#����xz���D�sv���**T½��-c�?��Y	@�DjS���1�a���`�
�&J���8�z�����[��G-��� _���k���d�iG�5�\���K׎"cY�]!�� I�S�U,
�h�C��ȃf�7���k!T|� �3��;�����Њ��v�j��������R�����h�-G���=!G��@�d�1ѵ�g�mNx311���޸�>Z�:zT��:�]�ȋ6-�h$��cx�&����N�h棟����r�-DR�8VP��J�����$��S�P���Mo�M2ȅ@�G�P!9�!�&��DO3ð?������Lٞr��v�T�5�l�GK��nq���\ˢ���B�0K{P�0�9�wrt����h�=�,P�)kgUzj��-�@���c.�(�9�_j��E:��s���4�v�0����ֺ�X��Ø3�+��`Y�S��̿�F��u�=`���1���a�7��.}9��WC;�?n��V_٘+��l~������?!� �H���j)��q굡w�� C�gZ<\KN����������Ό��
/��ۏ%&-n���B��+M{�sӇR�o�@���1��[�<$t�1�5���=_l�~��n�W��Е#���6.�mb��[1��I~��b�~�ͨ쎾ZK���so�&�4�D�D�v׃�p�#����P<	�����~�'ha���O�͙�z���{�Nת�Z=�D�����ol�1˝�iW��]��MKFD� F�o��)��q����|�33l��M�u�a���)Ô]����7�d�f�����G>�h���Z������$�^T(Z &*����.�̷���N����ơ�
�b-��ߓ�v�O��Qd��b߭�^����Cn��@~���Ac����6>Q=�B�y+�MC۞������A���RK&�pS�K�g`:��#����#H���a+��Nt"�p�q�o<�܌�6��R�!I�n \.H6�vz��?��?V��OX�Q�`�6�'~�ޗ�0s_}�~f�c^�)U��0�y�@'��n�W�� ��I�OÍ|n�8��m]@�)�C�3�\-�F�4�gx�
1����Ί�Z�}������)�J@ȝˮ�ݫ�#-�[*��`���dɹDI+��`��Yb���]��Ք���nX>�PK   ��X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   ��XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ��X�l�b�  �,     jsons/user_defined.json�Y�n�H�A��&�~�bev=_��F�A0�&�c2�PT�F�ߢ.�ؼ��1f���$Q�b�N���q�0����r�?2��g��7_-�?p�GKל���c����7���G��d��ֵ�Fg岨����KY=�%���Ɵ�V��;����h��ױ�Hpi���* *�BLr��
.X�$3�Ώ�_�U>��N�_�i�%�
\Ĕ�Ǟ!�A2x���*�p2/��uyZ�p��`��T��f�B"��0c��ls�</N�P������4_�g�ᤜAtƔ$�6p��{��	gF�5�:��"������c]��47T۪�,ys�g�lMe�q���`p�/����hƸxr^���]Y���q]-!�3�|s�<�v��u�p��1W{|yr�g6y�����ϫ]����f�̃��yU�}U�D�d�b�-D|����Ib;[6�(�~��՛\�+�_'����t����"o�l�U��2��<m���Ϝ-����������X�e�_�6�#�K ��o��$�{��(�ik"����Ԧw~�D߈�F�7���uzܬ��7/��|Y��e���3d��HgGF{��T��2�bɉ�%#x&�8�(��@����ͳ�E%
>��3�H�Lg�B+�|�8�S��0U��9�.[O���
=�ɟO�I�
]q�U��L�wU!�a��)��'6�l��y=:-�es��*d۩���o�i���ix2(��̤�ҭ*�C?P��G�������ʿ��Ue>���H(k���ʐ5�@�c>�X�Z�V8C�:���LbPU2ku�!��40̔s@j!-��sdi�(,dP���Eh)d���N-����6̟Ќ��K�ɑ�,��<�����a���s!��{h������	吖GDA(7{�	��g-x�IB�4�_��^xނWT'X(�c�E��{��-1�@�cXB�t�Y�9dAj(ؚ�}�X�T�`�d��RM*��z>A��]��^C�eH�I�1�iK��]�2-C�I��(���Qx(z��_��o�� 5_!�@#��#mj�o����㭾��W��6�	^�J�h��qjӛ��v��� �N�ڂ�X� �`9[?k���OA���]6�?�w�Ɩ﫞����Z�dn��zU��~[�Ɩ���ml�`�;���,�ѿOЪ%�3QO��W��Ge]�A�äU�f�Q�H����mLg�p��h��Lg�P�,��f��DpLg4�̴�ǜ�XrD<�9�Ns������Rl�!��^��l(��Er��_�D*,[��S�ߞ�2���Y��G��3@#\�7�����HW���~9;-���/~tvy#��O���ǹ��*����W��O3$t�eJ�,Z�#�{���!�AVgq�1��:&iD�C�D����(���I.����J$�B��#�tI�oB<,��E$�Ǔ��珺?�@���#<���=��۝�#<����@p�m�#<Y��].L����|�5���rz~[Wv�#=h�4eڃd�!�,Ao^�&��[��;���]�&U�̋rts~�L���*���*g�=��(˜��!%���Sd1u �P��%�il]
4��TP_�-2(S�K�r貭�������c��:^垂EM"���j�q�3����o�o>��/!"̻a������_�^{��>Hp�`Y��7y[�z�vPGa���U��ˠ�JCq�-���Q:�/����a�s̃vy4.�'��h\�O6QmJѸܟ,�ڄ�q�?�l���{A����M�����o$v2T I�V�������EX�$W�[����>�-�OZ�59�����!Z*���vh��D���m���v��Gms��HTُڦ�JbP����-��_i�p�H�~z������b�%#Q���:�KE�⾁c7`��I�E�q�rL;��]��c��/٩N�	i�������A�uv��oz>��PK   ��X��OZ%  j            ��    cirkitFile.jsonPK   ��X�<1	}�  � /           ��R  images/02d8db12-ba28-4e49-8e56-db179b980a39.pngPK   ��XWC��)�  � /           ��� images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK   ��Xx�آ  �  /           ���� images/0fa89018-bbd7-413a-af56-bcf37033748d.pngPK   ��X��_8
  3
  /           ���� images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK   ��X��MY��  �  /           ��� images/6e704699-d8e8-4ba8-9ba1-d4b639f353b6.pngPK   ��X(	��I�  &�  /           ��Nv images/9311ee57-74f3-4b31-a8d5-48402682b362.pngPK   ��X`$} [ /           ��� images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK   ��X�w3.  )  /           ��J�	 images/b3ba8064-1e10-4daf-8b84-7882f41f3c09.pngPK   ��X$7h�!  �!  /           ��Ŧ	 images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK   ��XKm���[ � /           ���	 images/e677f489-379d-40e3-bb59-6fe87b8e7dd0.pngPK   ��X�+�s;  z;  /           �� % images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK   ��XP��/�  ǽ  /           ���` images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK   ��X�l�b�  �,             ��> jsons/user_defined.jsonPK      �  T   